`timescale 1ns / 1ps

// show pixel(x, y) on the screen
module graphic(
    input wire  clk, reset,
    input wire  [10:0] x, y,
    input wire  BtnL,
    input wire  BtnR,
    input wire  BtnU,
    input wire  BtnD,
    output wire [7:0]  rgb
);

    // colors: [B1 B2 G1 G2 G3 R1 R2 R3]
    localparam COLOR_BG   = 8'b01001000;
    localparam COLOR_LINE = 8'b11100001;
    localparam COLOR_LARROW = 8'b11011101;
    localparam COLOR_RARROW = 8'b10010111;
    localparam COLOR_UARROW = 8'b00101011;
    localparam COLOR_DARROW = 8'b1011011;
    localparam COLOR_NULL = 8'b00000000;
    

    localparam U_BOUND = 11'd40;
    localparam D_BOUND = 11'd440;
    localparam H_ARR_W = 11'd40;
    localparam H_ARR_H = 11'd10;
    localparam V_ARR_W = 11'd10;
    localparam V_ARR_H = 11'd40;
    localparam U_ARR_X = 11'd128;
    localparam D_ARR_X = 11'd256;
    localparam L_ARR_X = 11'd384;
    localparam R_ARR_X = 11'd512;
    localparam SCORE_LINE_WIDTH = 11'd2;
    localparam SCORE_LINE_Y = 11'd440;

    localparam ARR_V = 10'd1;
    localparam SCORE_TOLERANCE = 11'd5;

    localparam MAX_ARROWS = 32;
    reg [10:0] score;
    reg [10:0] UArrows [MAX_ARROWS - 1:0];
    reg [10:0] LArrows [MAX_ARROWS - 1:0];
    reg [10:0] DArrows [MAX_ARROWS - 1:0];
    reg [10:0] RArrows [MAX_ARROWS - 1:0];
    reg [4:0] Uloc, Dloc, Lloc, Rloc;
    integer i;

    wire nclk;
    wire nclkedge;
    note_clk nclkgen(.clk(clk), .out_clk(nclk));
    edgedetect nced(.clk(clk), .sig(nclk), .possig(nclkedge));

    wire [4:0] rand;
    lfsr randgen(.clk(clk), .rst_n(reset));

    reg [7:0] rgb_now;
    wire clk_frame = (x == 0 && y == 0);
    always @(posedge clk) begin
        rand = rand + 1;

        if (reset) begin
            for (i = 0; i < MAX_ARROWS; i = i+1) begin
                UArrows[i] = 0;
                LArrows[i] = 0;
                DArrows[i] = 0;
                RArrows[i] = 0;
            end
            Uloc = 0;
            Dloc = 0;
            Lloc = 0;
            Rloc = 0;
            score = 0;
        end

        if (clk_frame) begin

            //generate new arrow every at certain frequency randomly choose which arrow type
            if(nclkedge) begin
                case rand[1:0]
                    0: begin
                        UArrows[Uloc] = U_BOUND;
                        Uloc = Uloc + 1;
                    end
                    1: begin
                        DArrows[Dloc] = U_BOUND;
                        Dloc = Dloc + 1;
                    end
                    2: begin
                        RArrows[Rloc] = U_BOUND;
                        Rloc = Rloc + 1;
                    end
                    3: begin
                        LArrows[Lloc] = U_BOUND;
                        Lloc = Lloc + 1;
                    end
                endcase
            end

            //check for correct presses
            for (i = 0; i < MAX_ARROWS; i = i+1) begin
                if (BtnU && (UArrows[i] >= SCORE_LINE_Y - SCORE_TOLERANCE && UArrows[i] <= SCORE_LINE_Y + SCORE_TOLERANCE)) begin
                    UArrows[i] = 0;
                    score = score + 1;
                end
                if (BtnD && (DArrows[i] >= SCORE_LINE_Y - SCORE_TOLERANCE && DArrows[i] <= SCORE_LINE_Y + SCORE_TOLERANCE)) begin
                    DArrows[i] = 0;
                    score = score + 1;
                end
                if (BtnL && (LArrows[i] >= SCORE_LINE_Y - SCORE_TOLERANCE && LArrows[i] <= SCORE_LINE_Y + SCORE_TOLERANCE)) begin
                    LArrows[i] = 0;
                    score = score + 1;
                end
                if (BtnR && (RArrows[i] >= SCORE_LINE_Y - SCORE_TOLERANCE && RArrows[i] <= SCORE_LINE_Y + SCORE_TOLERANCE)) begin
                    RArrows[i] = 0;
                    score = score + 1;
                end
            end


            //move arrows down
            for (i = 0; i < MAX_ARROWS; i = i+1) begin
                if (UArrows[i] != 0) begin
                    UArrows[i] = UArrows[i] + ARR_V;
                end
                if (DArrows[i] != 0) begin
                    DArrows[i] = DArrows[i] + ARR_V;
                end
                if (RArrows[i] != 0) begin
                    RArrows[i] = RArrows[i] + ARR_V;
                end
                if (LArrows[i] != 0) begin
                    LArrows[i] = LArrows[i] + ARR_V;
                end
            end
        end

        if (x >= 0 && y >= 0 && x < 640 && y < 480) begin

            rgb_now <= COLOR_BG;

            //arrows
            for (i = 0; i < MAX_ARROWS; i = i+1) begin
                if ((UArrows[i] != 0) && (x >= U_ARR_X - V_ARR_W/2 && x <= U_ARR_X + V_ARR_W/2) && (y >= UArrows[i] - V_ARR_H/2 && y <= UArrows[i] + V_ARR_H/2)) begin
                    rgb_now <= COLOR_UARROW;
                end
                if ((DArrows[i] != 0) && (x >= D_ARR_X - V_ARR_W/2 && x <= D_ARR_X + V_ARR_W/2) && (y >= DArrows[i] - V_ARR_H/2 && y <= DArrows[i] + V_ARR_H/2)) begin
                    rgb_now <= COLOR_DARROW;
                end
                if ((LArrows[i] != 0) && (x >= L_ARR_X - H_ARR_W/2 && x <= L_ARR_X + H_ARR_W/2) && (y >= LArrows[i] - H_ARR_H/2 && y <= LArrows[i] + H_ARR_H/2)) begin
                    rgb_now <= COLOR_LARROW;
                end
                if ((UArrows[i] != 0) && (x >= R_ARR_X - H_ARR_W/2 && x <= R_ARR_X + H_ARR_W/2) && (y >= RArrows[i] - H_ARR_H/2 && y <= RArrows[i] + H_ARR_H/2)) begin
                    rgb_now <= COLOR_RARROW;
                end
            end

            //score line
            if (y >= SCORE_LINE_Y - SCORE_LINE_WIDTH/2 && y <= SCORE_LINE_Y + SCORE_LINE_WIDTH/2) begin
                rgb_now <= COLOR_LINE;
            end

        end else begin
            // outside of the display area, fill black
            rgb_now <= COLOR_NULL;
        end
    end

    assign rgb = rgb_now;

endmodule