`timescale 1ns / 1ps

module BtoBCD(
    input clk, [15:0] bin,
    output reg [15:0] bcd
    );
    always @(posedge clk) begin
        case(bin)
            1: bcd <= 16'h0001;
            2: bcd <= 16'h0002;
            3: bcd <= 16'h0003;
            4: bcd <= 16'h0004;
            5: bcd <= 16'h0005;
            6: bcd <= 16'h0006;
            7: bcd <= 16'h0007;
            8: bcd <= 16'h0008;
            9: bcd <= 16'h0009;
            10: bcd <= 16'h0010;
            11: bcd <= 16'h0011;
            12: bcd <= 16'h0012;
            13: bcd <= 16'h0013;
            14: bcd <= 16'h0014;
            15: bcd <= 16'h0015;
            16: bcd <= 16'h0016;
            17: bcd <= 16'h0017;
            18: bcd <= 16'h0018;
            19: bcd <= 16'h0019;
            20: bcd <= 16'h0020;
            21: bcd <= 16'h0021;
            22: bcd <= 16'h0022;
            23: bcd <= 16'h0023;
            24: bcd <= 16'h0024;
            25: bcd <= 16'h0025;
            26: bcd <= 16'h0026;
            27: bcd <= 16'h0027;
            28: bcd <= 16'h0028;
            29: bcd <= 16'h0029;
            30: bcd <= 16'h0030;
            31: bcd <= 16'h0031;
            32: bcd <= 16'h0032;
            33: bcd <= 16'h0033;
            34: bcd <= 16'h0034;
            35: bcd <= 16'h0035;
            36: bcd <= 16'h0036;
            37: bcd <= 16'h0037;
            38: bcd <= 16'h0038;
            39: bcd <= 16'h0039;
            40: bcd <= 16'h0040;
            41: bcd <= 16'h0041;
            42: bcd <= 16'h0042;
            43: bcd <= 16'h0043;
            44: bcd <= 16'h0044;
            45: bcd <= 16'h0045;
            46: bcd <= 16'h0046;
            47: bcd <= 16'h0047;
            48: bcd <= 16'h0048;
            49: bcd <= 16'h0049;
            50: bcd <= 16'h0050;
            51: bcd <= 16'h0051;
            52: bcd <= 16'h0052;
            53: bcd <= 16'h0053;
            54: bcd <= 16'h0054;
            55: bcd <= 16'h0055;
            56: bcd <= 16'h0056;
            57: bcd <= 16'h0057;
            58: bcd <= 16'h0058;
            59: bcd <= 16'h0059;
            60: bcd <= 16'h0060;
            61: bcd <= 16'h0061;
            62: bcd <= 16'h0062;
            63: bcd <= 16'h0063;
            64: bcd <= 16'h0064;
            65: bcd <= 16'h0065;
            66: bcd <= 16'h0066;
            67: bcd <= 16'h0067;
            68: bcd <= 16'h0068;
            69: bcd <= 16'h0069;
            70: bcd <= 16'h0070;
            71: bcd <= 16'h0071;
            72: bcd <= 16'h0072;
            73: bcd <= 16'h0073;
            74: bcd <= 16'h0074;
            75: bcd <= 16'h0075;
            76: bcd <= 16'h0076;
            77: bcd <= 16'h0077;
            78: bcd <= 16'h0078;
            79: bcd <= 16'h0079;
            80: bcd <= 16'h0080;
            81: bcd <= 16'h0081;
            82: bcd <= 16'h0082;
            83: bcd <= 16'h0083;
            84: bcd <= 16'h0084;
            85: bcd <= 16'h0085;
            86: bcd <= 16'h0086;
            87: bcd <= 16'h0087;
            88: bcd <= 16'h0088;
            89: bcd <= 16'h0089;
            90: bcd <= 16'h0090;
            91: bcd <= 16'h0091;
            92: bcd <= 16'h0092;
            93: bcd <= 16'h0093;
            94: bcd <= 16'h0094;
            95: bcd <= 16'h0095;
            96: bcd <= 16'h0096;
            97: bcd <= 16'h0097;
            98: bcd <= 16'h0098;
            99: bcd <= 16'h0099;
            100: bcd <= 16'h0100;
            101: bcd <= 16'h0101;
            102: bcd <= 16'h0102;
            103: bcd <= 16'h0103;
            104: bcd <= 16'h0104;
            105: bcd <= 16'h0105;
            106: bcd <= 16'h0106;
            107: bcd <= 16'h0107;
            108: bcd <= 16'h0108;
            109: bcd <= 16'h0109;
            110: bcd <= 16'h0110;
            111: bcd <= 16'h0111;
            112: bcd <= 16'h0112;
            113: bcd <= 16'h0113;
            114: bcd <= 16'h0114;
            115: bcd <= 16'h0115;
            116: bcd <= 16'h0116;
            117: bcd <= 16'h0117;
            118: bcd <= 16'h0118;
            119: bcd <= 16'h0119;
            120: bcd <= 16'h0120;
            121: bcd <= 16'h0121;
            122: bcd <= 16'h0122;
            123: bcd <= 16'h0123;
            124: bcd <= 16'h0124;
            125: bcd <= 16'h0125;
            126: bcd <= 16'h0126;
            127: bcd <= 16'h0127;
            128: bcd <= 16'h0128;
            129: bcd <= 16'h0129;
            130: bcd <= 16'h0130;
            131: bcd <= 16'h0131;
            132: bcd <= 16'h0132;
            133: bcd <= 16'h0133;
            134: bcd <= 16'h0134;
            135: bcd <= 16'h0135;
            136: bcd <= 16'h0136;
            137: bcd <= 16'h0137;
            138: bcd <= 16'h0138;
            139: bcd <= 16'h0139;
            140: bcd <= 16'h0140;
            141: bcd <= 16'h0141;
            142: bcd <= 16'h0142;
            143: bcd <= 16'h0143;
            144: bcd <= 16'h0144;
            145: bcd <= 16'h0145;
            146: bcd <= 16'h0146;
            147: bcd <= 16'h0147;
            148: bcd <= 16'h0148;
            149: bcd <= 16'h0149;
            150: bcd <= 16'h0150;
            151: bcd <= 16'h0151;
            152: bcd <= 16'h0152;
            153: bcd <= 16'h0153;
            154: bcd <= 16'h0154;
            155: bcd <= 16'h0155;
            156: bcd <= 16'h0156;
            157: bcd <= 16'h0157;
            158: bcd <= 16'h0158;
            159: bcd <= 16'h0159;
            160: bcd <= 16'h0160;
            161: bcd <= 16'h0161;
            162: bcd <= 16'h0162;
            163: bcd <= 16'h0163;
            164: bcd <= 16'h0164;
            165: bcd <= 16'h0165;
            166: bcd <= 16'h0166;
            167: bcd <= 16'h0167;
            168: bcd <= 16'h0168;
            169: bcd <= 16'h0169;
            170: bcd <= 16'h0170;
            171: bcd <= 16'h0171;
            172: bcd <= 16'h0172;
            173: bcd <= 16'h0173;
            174: bcd <= 16'h0174;
            175: bcd <= 16'h0175;
            176: bcd <= 16'h0176;
            177: bcd <= 16'h0177;
            178: bcd <= 16'h0178;
            179: bcd <= 16'h0179;
            180: bcd <= 16'h0180;
            181: bcd <= 16'h0181;
            182: bcd <= 16'h0182;
            183: bcd <= 16'h0183;
            184: bcd <= 16'h0184;
            185: bcd <= 16'h0185;
            186: bcd <= 16'h0186;
            187: bcd <= 16'h0187;
            188: bcd <= 16'h0188;
            189: bcd <= 16'h0189;
            190: bcd <= 16'h0190;
            191: bcd <= 16'h0191;
            192: bcd <= 16'h0192;
            193: bcd <= 16'h0193;
            194: bcd <= 16'h0194;
            195: bcd <= 16'h0195;
            196: bcd <= 16'h0196;
            197: bcd <= 16'h0197;
            198: bcd <= 16'h0198;
            199: bcd <= 16'h0199;
            200: bcd <= 16'h0200;
            201: bcd <= 16'h0201;
            202: bcd <= 16'h0202;
            203: bcd <= 16'h0203;
            204: bcd <= 16'h0204;
            205: bcd <= 16'h0205;
            206: bcd <= 16'h0206;
            207: bcd <= 16'h0207;
            208: bcd <= 16'h0208;
            209: bcd <= 16'h0209;
            210: bcd <= 16'h0210;
            211: bcd <= 16'h0211;
            212: bcd <= 16'h0212;
            213: bcd <= 16'h0213;
            214: bcd <= 16'h0214;
            215: bcd <= 16'h0215;
            216: bcd <= 16'h0216;
            217: bcd <= 16'h0217;
            218: bcd <= 16'h0218;
            219: bcd <= 16'h0219;
            220: bcd <= 16'h0220;
            221: bcd <= 16'h0221;
            222: bcd <= 16'h0222;
            223: bcd <= 16'h0223;
            224: bcd <= 16'h0224;
            225: bcd <= 16'h0225;
            226: bcd <= 16'h0226;
            227: bcd <= 16'h0227;
            228: bcd <= 16'h0228;
            229: bcd <= 16'h0229;
            230: bcd <= 16'h0230;
            231: bcd <= 16'h0231;
            232: bcd <= 16'h0232;
            233: bcd <= 16'h0233;
            234: bcd <= 16'h0234;
            235: bcd <= 16'h0235;
            236: bcd <= 16'h0236;
            237: bcd <= 16'h0237;
            238: bcd <= 16'h0238;
            239: bcd <= 16'h0239;
            240: bcd <= 16'h0240;
            241: bcd <= 16'h0241;
            242: bcd <= 16'h0242;
            243: bcd <= 16'h0243;
            244: bcd <= 16'h0244;
            245: bcd <= 16'h0245;
            246: bcd <= 16'h0246;
            247: bcd <= 16'h0247;
            248: bcd <= 16'h0248;
            249: bcd <= 16'h0249;
            250: bcd <= 16'h0250;
            251: bcd <= 16'h0251;
            252: bcd <= 16'h0252;
            253: bcd <= 16'h0253;
            254: bcd <= 16'h0254;
            255: bcd <= 16'h0255;
            256: bcd <= 16'h0256;
            257: bcd <= 16'h0257;
            258: bcd <= 16'h0258;
            259: bcd <= 16'h0259;
            260: bcd <= 16'h0260;
            261: bcd <= 16'h0261;
            262: bcd <= 16'h0262;
            263: bcd <= 16'h0263;
            264: bcd <= 16'h0264;
            265: bcd <= 16'h0265;
            266: bcd <= 16'h0266;
            267: bcd <= 16'h0267;
            268: bcd <= 16'h0268;
            269: bcd <= 16'h0269;
            270: bcd <= 16'h0270;
            271: bcd <= 16'h0271;
            272: bcd <= 16'h0272;
            273: bcd <= 16'h0273;
            274: bcd <= 16'h0274;
            275: bcd <= 16'h0275;
            276: bcd <= 16'h0276;
            277: bcd <= 16'h0277;
            278: bcd <= 16'h0278;
            279: bcd <= 16'h0279;
            280: bcd <= 16'h0280;
            281: bcd <= 16'h0281;
            282: bcd <= 16'h0282;
            283: bcd <= 16'h0283;
            284: bcd <= 16'h0284;
            285: bcd <= 16'h0285;
            286: bcd <= 16'h0286;
            287: bcd <= 16'h0287;
            288: bcd <= 16'h0288;
            289: bcd <= 16'h0289;
            290: bcd <= 16'h0290;
            291: bcd <= 16'h0291;
            292: bcd <= 16'h0292;
            293: bcd <= 16'h0293;
            294: bcd <= 16'h0294;
            295: bcd <= 16'h0295;
            296: bcd <= 16'h0296;
            297: bcd <= 16'h0297;
            298: bcd <= 16'h0298;
            299: bcd <= 16'h0299;
            300: bcd <= 16'h0300;
            301: bcd <= 16'h0301;
            302: bcd <= 16'h0302;
            303: bcd <= 16'h0303;
            304: bcd <= 16'h0304;
            305: bcd <= 16'h0305;
            306: bcd <= 16'h0306;
            307: bcd <= 16'h0307;
            308: bcd <= 16'h0308;
            309: bcd <= 16'h0309;
            310: bcd <= 16'h0310;
            311: bcd <= 16'h0311;
            312: bcd <= 16'h0312;
            313: bcd <= 16'h0313;
            314: bcd <= 16'h0314;
            315: bcd <= 16'h0315;
            316: bcd <= 16'h0316;
            317: bcd <= 16'h0317;
            318: bcd <= 16'h0318;
            319: bcd <= 16'h0319;
            320: bcd <= 16'h0320;
            321: bcd <= 16'h0321;
            322: bcd <= 16'h0322;
            323: bcd <= 16'h0323;
            324: bcd <= 16'h0324;
            325: bcd <= 16'h0325;
            326: bcd <= 16'h0326;
            327: bcd <= 16'h0327;
            328: bcd <= 16'h0328;
            329: bcd <= 16'h0329;
            330: bcd <= 16'h0330;
            331: bcd <= 16'h0331;
            332: bcd <= 16'h0332;
            333: bcd <= 16'h0333;
            334: bcd <= 16'h0334;
            335: bcd <= 16'h0335;
            336: bcd <= 16'h0336;
            337: bcd <= 16'h0337;
            338: bcd <= 16'h0338;
            339: bcd <= 16'h0339;
            340: bcd <= 16'h0340;
            341: bcd <= 16'h0341;
            342: bcd <= 16'h0342;
            343: bcd <= 16'h0343;
            344: bcd <= 16'h0344;
            345: bcd <= 16'h0345;
            346: bcd <= 16'h0346;
            347: bcd <= 16'h0347;
            348: bcd <= 16'h0348;
            349: bcd <= 16'h0349;
            350: bcd <= 16'h0350;
            351: bcd <= 16'h0351;
            352: bcd <= 16'h0352;
            353: bcd <= 16'h0353;
            354: bcd <= 16'h0354;
            355: bcd <= 16'h0355;
            356: bcd <= 16'h0356;
            357: bcd <= 16'h0357;
            358: bcd <= 16'h0358;
            359: bcd <= 16'h0359;
            360: bcd <= 16'h0360;
            361: bcd <= 16'h0361;
            362: bcd <= 16'h0362;
            363: bcd <= 16'h0363;
            364: bcd <= 16'h0364;
            365: bcd <= 16'h0365;
            366: bcd <= 16'h0366;
            367: bcd <= 16'h0367;
            368: bcd <= 16'h0368;
            369: bcd <= 16'h0369;
            370: bcd <= 16'h0370;
            371: bcd <= 16'h0371;
            372: bcd <= 16'h0372;
            373: bcd <= 16'h0373;
            374: bcd <= 16'h0374;
            375: bcd <= 16'h0375;
            376: bcd <= 16'h0376;
            377: bcd <= 16'h0377;
            378: bcd <= 16'h0378;
            379: bcd <= 16'h0379;
            380: bcd <= 16'h0380;
            381: bcd <= 16'h0381;
            382: bcd <= 16'h0382;
            383: bcd <= 16'h0383;
            384: bcd <= 16'h0384;
            385: bcd <= 16'h0385;
            386: bcd <= 16'h0386;
            387: bcd <= 16'h0387;
            388: bcd <= 16'h0388;
            389: bcd <= 16'h0389;
            390: bcd <= 16'h0390;
            391: bcd <= 16'h0391;
            392: bcd <= 16'h0392;
            393: bcd <= 16'h0393;
            394: bcd <= 16'h0394;
            395: bcd <= 16'h0395;
            396: bcd <= 16'h0396;
            397: bcd <= 16'h0397;
            398: bcd <= 16'h0398;
            399: bcd <= 16'h0399;
            400: bcd <= 16'h0400;
            401: bcd <= 16'h0401;
            402: bcd <= 16'h0402;
            403: bcd <= 16'h0403;
            404: bcd <= 16'h0404;
            405: bcd <= 16'h0405;
            406: bcd <= 16'h0406;
            407: bcd <= 16'h0407;
            408: bcd <= 16'h0408;
            409: bcd <= 16'h0409;
            410: bcd <= 16'h0410;
            411: bcd <= 16'h0411;
            412: bcd <= 16'h0412;
            413: bcd <= 16'h0413;
            414: bcd <= 16'h0414;
            415: bcd <= 16'h0415;
            416: bcd <= 16'h0416;
            417: bcd <= 16'h0417;
            418: bcd <= 16'h0418;
            419: bcd <= 16'h0419;
            420: bcd <= 16'h0420;
            421: bcd <= 16'h0421;
            422: bcd <= 16'h0422;
            423: bcd <= 16'h0423;
            424: bcd <= 16'h0424;
            425: bcd <= 16'h0425;
            426: bcd <= 16'h0426;
            427: bcd <= 16'h0427;
            428: bcd <= 16'h0428;
            429: bcd <= 16'h0429;
            430: bcd <= 16'h0430;
            431: bcd <= 16'h0431;
            432: bcd <= 16'h0432;
            433: bcd <= 16'h0433;
            434: bcd <= 16'h0434;
            435: bcd <= 16'h0435;
            436: bcd <= 16'h0436;
            437: bcd <= 16'h0437;
            438: bcd <= 16'h0438;
            439: bcd <= 16'h0439;
            440: bcd <= 16'h0440;
            441: bcd <= 16'h0441;
            442: bcd <= 16'h0442;
            443: bcd <= 16'h0443;
            444: bcd <= 16'h0444;
            445: bcd <= 16'h0445;
            446: bcd <= 16'h0446;
            447: bcd <= 16'h0447;
            448: bcd <= 16'h0448;
            449: bcd <= 16'h0449;
            450: bcd <= 16'h0450;
            451: bcd <= 16'h0451;
            452: bcd <= 16'h0452;
            453: bcd <= 16'h0453;
            454: bcd <= 16'h0454;
            455: bcd <= 16'h0455;
            456: bcd <= 16'h0456;
            457: bcd <= 16'h0457;
            458: bcd <= 16'h0458;
            459: bcd <= 16'h0459;
            460: bcd <= 16'h0460;
            461: bcd <= 16'h0461;
            462: bcd <= 16'h0462;
            463: bcd <= 16'h0463;
            464: bcd <= 16'h0464;
            465: bcd <= 16'h0465;
            466: bcd <= 16'h0466;
            467: bcd <= 16'h0467;
            468: bcd <= 16'h0468;
            469: bcd <= 16'h0469;
            470: bcd <= 16'h0470;
            471: bcd <= 16'h0471;
            472: bcd <= 16'h0472;
            473: bcd <= 16'h0473;
            474: bcd <= 16'h0474;
            475: bcd <= 16'h0475;
            476: bcd <= 16'h0476;
            477: bcd <= 16'h0477;
            478: bcd <= 16'h0478;
            479: bcd <= 16'h0479;
            480: bcd <= 16'h0480;
            481: bcd <= 16'h0481;
            482: bcd <= 16'h0482;
            483: bcd <= 16'h0483;
            484: bcd <= 16'h0484;
            485: bcd <= 16'h0485;
            486: bcd <= 16'h0486;
            487: bcd <= 16'h0487;
            488: bcd <= 16'h0488;
            489: bcd <= 16'h0489;
            490: bcd <= 16'h0490;
            491: bcd <= 16'h0491;
            492: bcd <= 16'h0492;
            493: bcd <= 16'h0493;
            494: bcd <= 16'h0494;
            495: bcd <= 16'h0495;
            496: bcd <= 16'h0496;
            497: bcd <= 16'h0497;
            498: bcd <= 16'h0498;
            499: bcd <= 16'h0499;
            500: bcd <= 16'h0500;
            501: bcd <= 16'h0501;
            502: bcd <= 16'h0502;
            503: bcd <= 16'h0503;
            504: bcd <= 16'h0504;
            505: bcd <= 16'h0505;
            506: bcd <= 16'h0506;
            507: bcd <= 16'h0507;
            508: bcd <= 16'h0508;
            509: bcd <= 16'h0509;
            510: bcd <= 16'h0510;
            511: bcd <= 16'h0511;
            512: bcd <= 16'h0512;
            513: bcd <= 16'h0513;
            514: bcd <= 16'h0514;
            515: bcd <= 16'h0515;
            516: bcd <= 16'h0516;
            517: bcd <= 16'h0517;
            518: bcd <= 16'h0518;
            519: bcd <= 16'h0519;
            520: bcd <= 16'h0520;
            521: bcd <= 16'h0521;
            522: bcd <= 16'h0522;
            523: bcd <= 16'h0523;
            524: bcd <= 16'h0524;
            525: bcd <= 16'h0525;
            526: bcd <= 16'h0526;
            527: bcd <= 16'h0527;
            528: bcd <= 16'h0528;
            529: bcd <= 16'h0529;
            530: bcd <= 16'h0530;
            531: bcd <= 16'h0531;
            532: bcd <= 16'h0532;
            533: bcd <= 16'h0533;
            534: bcd <= 16'h0534;
            535: bcd <= 16'h0535;
            536: bcd <= 16'h0536;
            537: bcd <= 16'h0537;
            538: bcd <= 16'h0538;
            539: bcd <= 16'h0539;
            540: bcd <= 16'h0540;
            541: bcd <= 16'h0541;
            542: bcd <= 16'h0542;
            543: bcd <= 16'h0543;
            544: bcd <= 16'h0544;
            545: bcd <= 16'h0545;
            546: bcd <= 16'h0546;
            547: bcd <= 16'h0547;
            548: bcd <= 16'h0548;
            549: bcd <= 16'h0549;
            550: bcd <= 16'h0550;
            551: bcd <= 16'h0551;
            552: bcd <= 16'h0552;
            553: bcd <= 16'h0553;
            554: bcd <= 16'h0554;
            555: bcd <= 16'h0555;
            556: bcd <= 16'h0556;
            557: bcd <= 16'h0557;
            558: bcd <= 16'h0558;
            559: bcd <= 16'h0559;
            560: bcd <= 16'h0560;
            561: bcd <= 16'h0561;
            562: bcd <= 16'h0562;
            563: bcd <= 16'h0563;
            564: bcd <= 16'h0564;
            565: bcd <= 16'h0565;
            566: bcd <= 16'h0566;
            567: bcd <= 16'h0567;
            568: bcd <= 16'h0568;
            569: bcd <= 16'h0569;
            570: bcd <= 16'h0570;
            571: bcd <= 16'h0571;
            572: bcd <= 16'h0572;
            573: bcd <= 16'h0573;
            574: bcd <= 16'h0574;
            575: bcd <= 16'h0575;
            576: bcd <= 16'h0576;
            577: bcd <= 16'h0577;
            578: bcd <= 16'h0578;
            579: bcd <= 16'h0579;
            580: bcd <= 16'h0580;
            581: bcd <= 16'h0581;
            582: bcd <= 16'h0582;
            583: bcd <= 16'h0583;
            584: bcd <= 16'h0584;
            585: bcd <= 16'h0585;
            586: bcd <= 16'h0586;
            587: bcd <= 16'h0587;
            588: bcd <= 16'h0588;
            589: bcd <= 16'h0589;
            590: bcd <= 16'h0590;
            591: bcd <= 16'h0591;
            592: bcd <= 16'h0592;
            593: bcd <= 16'h0593;
            594: bcd <= 16'h0594;
            595: bcd <= 16'h0595;
            596: bcd <= 16'h0596;
            597: bcd <= 16'h0597;
            598: bcd <= 16'h0598;
            599: bcd <= 16'h0599;
            600: bcd <= 16'h0600;
            601: bcd <= 16'h0601;
            602: bcd <= 16'h0602;
            603: bcd <= 16'h0603;
            604: bcd <= 16'h0604;
            605: bcd <= 16'h0605;
            606: bcd <= 16'h0606;
            607: bcd <= 16'h0607;
            608: bcd <= 16'h0608;
            609: bcd <= 16'h0609;
            610: bcd <= 16'h0610;
            611: bcd <= 16'h0611;
            612: bcd <= 16'h0612;
            613: bcd <= 16'h0613;
            614: bcd <= 16'h0614;
            615: bcd <= 16'h0615;
            616: bcd <= 16'h0616;
            617: bcd <= 16'h0617;
            618: bcd <= 16'h0618;
            619: bcd <= 16'h0619;
            620: bcd <= 16'h0620;
            621: bcd <= 16'h0621;
            622: bcd <= 16'h0622;
            623: bcd <= 16'h0623;
            624: bcd <= 16'h0624;
            625: bcd <= 16'h0625;
            626: bcd <= 16'h0626;
            627: bcd <= 16'h0627;
            628: bcd <= 16'h0628;
            629: bcd <= 16'h0629;
            630: bcd <= 16'h0630;
            631: bcd <= 16'h0631;
            632: bcd <= 16'h0632;
            633: bcd <= 16'h0633;
            634: bcd <= 16'h0634;
            635: bcd <= 16'h0635;
            636: bcd <= 16'h0636;
            637: bcd <= 16'h0637;
            638: bcd <= 16'h0638;
            639: bcd <= 16'h0639;
            640: bcd <= 16'h0640;
            641: bcd <= 16'h0641;
            642: bcd <= 16'h0642;
            643: bcd <= 16'h0643;
            644: bcd <= 16'h0644;
            645: bcd <= 16'h0645;
            646: bcd <= 16'h0646;
            647: bcd <= 16'h0647;
            648: bcd <= 16'h0648;
            649: bcd <= 16'h0649;
            650: bcd <= 16'h0650;
            651: bcd <= 16'h0651;
            652: bcd <= 16'h0652;
            653: bcd <= 16'h0653;
            654: bcd <= 16'h0654;
            655: bcd <= 16'h0655;
            656: bcd <= 16'h0656;
            657: bcd <= 16'h0657;
            658: bcd <= 16'h0658;
            659: bcd <= 16'h0659;
            660: bcd <= 16'h0660;
            661: bcd <= 16'h0661;
            662: bcd <= 16'h0662;
            663: bcd <= 16'h0663;
            664: bcd <= 16'h0664;
            665: bcd <= 16'h0665;
            666: bcd <= 16'h0666;
            667: bcd <= 16'h0667;
            668: bcd <= 16'h0668;
            669: bcd <= 16'h0669;
            670: bcd <= 16'h0670;
            671: bcd <= 16'h0671;
            672: bcd <= 16'h0672;
            673: bcd <= 16'h0673;
            674: bcd <= 16'h0674;
            675: bcd <= 16'h0675;
            676: bcd <= 16'h0676;
            677: bcd <= 16'h0677;
            678: bcd <= 16'h0678;
            679: bcd <= 16'h0679;
            680: bcd <= 16'h0680;
            681: bcd <= 16'h0681;
            682: bcd <= 16'h0682;
            683: bcd <= 16'h0683;
            684: bcd <= 16'h0684;
            685: bcd <= 16'h0685;
            686: bcd <= 16'h0686;
            687: bcd <= 16'h0687;
            688: bcd <= 16'h0688;
            689: bcd <= 16'h0689;
            690: bcd <= 16'h0690;
            691: bcd <= 16'h0691;
            692: bcd <= 16'h0692;
            693: bcd <= 16'h0693;
            694: bcd <= 16'h0694;
            695: bcd <= 16'h0695;
            696: bcd <= 16'h0696;
            697: bcd <= 16'h0697;
            698: bcd <= 16'h0698;
            699: bcd <= 16'h0699;
            700: bcd <= 16'h0700;
            701: bcd <= 16'h0701;
            702: bcd <= 16'h0702;
            703: bcd <= 16'h0703;
            704: bcd <= 16'h0704;
            705: bcd <= 16'h0705;
            706: bcd <= 16'h0706;
            707: bcd <= 16'h0707;
            708: bcd <= 16'h0708;
            709: bcd <= 16'h0709;
            710: bcd <= 16'h0710;
            711: bcd <= 16'h0711;
            712: bcd <= 16'h0712;
            713: bcd <= 16'h0713;
            714: bcd <= 16'h0714;
            715: bcd <= 16'h0715;
            716: bcd <= 16'h0716;
            717: bcd <= 16'h0717;
            718: bcd <= 16'h0718;
            719: bcd <= 16'h0719;
            720: bcd <= 16'h0720;
            721: bcd <= 16'h0721;
            722: bcd <= 16'h0722;
            723: bcd <= 16'h0723;
            724: bcd <= 16'h0724;
            725: bcd <= 16'h0725;
            726: bcd <= 16'h0726;
            727: bcd <= 16'h0727;
            728: bcd <= 16'h0728;
            729: bcd <= 16'h0729;
            730: bcd <= 16'h0730;
            731: bcd <= 16'h0731;
            732: bcd <= 16'h0732;
            733: bcd <= 16'h0733;
            734: bcd <= 16'h0734;
            735: bcd <= 16'h0735;
            736: bcd <= 16'h0736;
            737: bcd <= 16'h0737;
            738: bcd <= 16'h0738;
            739: bcd <= 16'h0739;
            740: bcd <= 16'h0740;
            741: bcd <= 16'h0741;
            742: bcd <= 16'h0742;
            743: bcd <= 16'h0743;
            744: bcd <= 16'h0744;
            745: bcd <= 16'h0745;
            746: bcd <= 16'h0746;
            747: bcd <= 16'h0747;
            748: bcd <= 16'h0748;
            749: bcd <= 16'h0749;
            750: bcd <= 16'h0750;
            751: bcd <= 16'h0751;
            752: bcd <= 16'h0752;
            753: bcd <= 16'h0753;
            754: bcd <= 16'h0754;
            755: bcd <= 16'h0755;
            756: bcd <= 16'h0756;
            757: bcd <= 16'h0757;
            758: bcd <= 16'h0758;
            759: bcd <= 16'h0759;
            760: bcd <= 16'h0760;
            761: bcd <= 16'h0761;
            762: bcd <= 16'h0762;
            763: bcd <= 16'h0763;
            764: bcd <= 16'h0764;
            765: bcd <= 16'h0765;
            766: bcd <= 16'h0766;
            767: bcd <= 16'h0767;
            768: bcd <= 16'h0768;
            769: bcd <= 16'h0769;
            770: bcd <= 16'h0770;
            771: bcd <= 16'h0771;
            772: bcd <= 16'h0772;
            773: bcd <= 16'h0773;
            774: bcd <= 16'h0774;
            775: bcd <= 16'h0775;
            776: bcd <= 16'h0776;
            777: bcd <= 16'h0777;
            778: bcd <= 16'h0778;
            779: bcd <= 16'h0779;
            780: bcd <= 16'h0780;
            781: bcd <= 16'h0781;
            782: bcd <= 16'h0782;
            783: bcd <= 16'h0783;
            784: bcd <= 16'h0784;
            785: bcd <= 16'h0785;
            786: bcd <= 16'h0786;
            787: bcd <= 16'h0787;
            788: bcd <= 16'h0788;
            789: bcd <= 16'h0789;
            790: bcd <= 16'h0790;
            791: bcd <= 16'h0791;
            792: bcd <= 16'h0792;
            793: bcd <= 16'h0793;
            794: bcd <= 16'h0794;
            795: bcd <= 16'h0795;
            796: bcd <= 16'h0796;
            797: bcd <= 16'h0797;
            798: bcd <= 16'h0798;
            799: bcd <= 16'h0799;
            800: bcd <= 16'h0800;
            801: bcd <= 16'h0801;
            802: bcd <= 16'h0802;
            803: bcd <= 16'h0803;
            804: bcd <= 16'h0804;
            805: bcd <= 16'h0805;
            806: bcd <= 16'h0806;
            807: bcd <= 16'h0807;
            808: bcd <= 16'h0808;
            809: bcd <= 16'h0809;
            810: bcd <= 16'h0810;
            811: bcd <= 16'h0811;
            812: bcd <= 16'h0812;
            813: bcd <= 16'h0813;
            814: bcd <= 16'h0814;
            815: bcd <= 16'h0815;
            816: bcd <= 16'h0816;
            817: bcd <= 16'h0817;
            818: bcd <= 16'h0818;
            819: bcd <= 16'h0819;
            820: bcd <= 16'h0820;
            821: bcd <= 16'h0821;
            822: bcd <= 16'h0822;
            823: bcd <= 16'h0823;
            824: bcd <= 16'h0824;
            825: bcd <= 16'h0825;
            826: bcd <= 16'h0826;
            827: bcd <= 16'h0827;
            828: bcd <= 16'h0828;
            829: bcd <= 16'h0829;
            830: bcd <= 16'h0830;
            831: bcd <= 16'h0831;
            832: bcd <= 16'h0832;
            833: bcd <= 16'h0833;
            834: bcd <= 16'h0834;
            835: bcd <= 16'h0835;
            836: bcd <= 16'h0836;
            837: bcd <= 16'h0837;
            838: bcd <= 16'h0838;
            839: bcd <= 16'h0839;
            840: bcd <= 16'h0840;
            841: bcd <= 16'h0841;
            842: bcd <= 16'h0842;
            843: bcd <= 16'h0843;
            844: bcd <= 16'h0844;
            845: bcd <= 16'h0845;
            846: bcd <= 16'h0846;
            847: bcd <= 16'h0847;
            848: bcd <= 16'h0848;
            849: bcd <= 16'h0849;
            850: bcd <= 16'h0850;
            851: bcd <= 16'h0851;
            852: bcd <= 16'h0852;
            853: bcd <= 16'h0853;
            854: bcd <= 16'h0854;
            855: bcd <= 16'h0855;
            856: bcd <= 16'h0856;
            857: bcd <= 16'h0857;
            858: bcd <= 16'h0858;
            859: bcd <= 16'h0859;
            860: bcd <= 16'h0860;
            861: bcd <= 16'h0861;
            862: bcd <= 16'h0862;
            863: bcd <= 16'h0863;
            864: bcd <= 16'h0864;
            865: bcd <= 16'h0865;
            866: bcd <= 16'h0866;
            867: bcd <= 16'h0867;
            868: bcd <= 16'h0868;
            869: bcd <= 16'h0869;
            870: bcd <= 16'h0870;
            871: bcd <= 16'h0871;
            872: bcd <= 16'h0872;
            873: bcd <= 16'h0873;
            874: bcd <= 16'h0874;
            875: bcd <= 16'h0875;
            876: bcd <= 16'h0876;
            877: bcd <= 16'h0877;
            878: bcd <= 16'h0878;
            879: bcd <= 16'h0879;
            880: bcd <= 16'h0880;
            881: bcd <= 16'h0881;
            882: bcd <= 16'h0882;
            883: bcd <= 16'h0883;
            884: bcd <= 16'h0884;
            885: bcd <= 16'h0885;
            886: bcd <= 16'h0886;
            887: bcd <= 16'h0887;
            888: bcd <= 16'h0888;
            889: bcd <= 16'h0889;
            890: bcd <= 16'h0890;
            891: bcd <= 16'h0891;
            892: bcd <= 16'h0892;
            893: bcd <= 16'h0893;
            894: bcd <= 16'h0894;
            895: bcd <= 16'h0895;
            896: bcd <= 16'h0896;
            897: bcd <= 16'h0897;
            898: bcd <= 16'h0898;
            899: bcd <= 16'h0899;
            900: bcd <= 16'h0900;
            901: bcd <= 16'h0901;
            902: bcd <= 16'h0902;
            903: bcd <= 16'h0903;
            904: bcd <= 16'h0904;
            905: bcd <= 16'h0905;
            906: bcd <= 16'h0906;
            907: bcd <= 16'h0907;
            908: bcd <= 16'h0908;
            909: bcd <= 16'h0909;
            910: bcd <= 16'h0910;
            911: bcd <= 16'h0911;
            912: bcd <= 16'h0912;
            913: bcd <= 16'h0913;
            914: bcd <= 16'h0914;
            915: bcd <= 16'h0915;
            916: bcd <= 16'h0916;
            917: bcd <= 16'h0917;
            918: bcd <= 16'h0918;
            919: bcd <= 16'h0919;
            920: bcd <= 16'h0920;
            921: bcd <= 16'h0921;
            922: bcd <= 16'h0922;
            923: bcd <= 16'h0923;
            924: bcd <= 16'h0924;
            925: bcd <= 16'h0925;
            926: bcd <= 16'h0926;
            927: bcd <= 16'h0927;
            928: bcd <= 16'h0928;
            929: bcd <= 16'h0929;
            930: bcd <= 16'h0930;
            931: bcd <= 16'h0931;
            932: bcd <= 16'h0932;
            933: bcd <= 16'h0933;
            934: bcd <= 16'h0934;
            935: bcd <= 16'h0935;
            936: bcd <= 16'h0936;
            937: bcd <= 16'h0937;
            938: bcd <= 16'h0938;
            939: bcd <= 16'h0939;
            940: bcd <= 16'h0940;
            941: bcd <= 16'h0941;
            942: bcd <= 16'h0942;
            943: bcd <= 16'h0943;
            944: bcd <= 16'h0944;
            945: bcd <= 16'h0945;
            946: bcd <= 16'h0946;
            947: bcd <= 16'h0947;
            948: bcd <= 16'h0948;
            949: bcd <= 16'h0949;
            950: bcd <= 16'h0950;
            951: bcd <= 16'h0951;
            952: bcd <= 16'h0952;
            953: bcd <= 16'h0953;
            954: bcd <= 16'h0954;
            955: bcd <= 16'h0955;
            956: bcd <= 16'h0956;
            957: bcd <= 16'h0957;
            958: bcd <= 16'h0958;
            959: bcd <= 16'h0959;
            960: bcd <= 16'h0960;
            961: bcd <= 16'h0961;
            962: bcd <= 16'h0962;
            963: bcd <= 16'h0963;
            964: bcd <= 16'h0964;
            965: bcd <= 16'h0965;
            966: bcd <= 16'h0966;
            967: bcd <= 16'h0967;
            968: bcd <= 16'h0968;
            969: bcd <= 16'h0969;
            970: bcd <= 16'h0970;
            971: bcd <= 16'h0971;
            972: bcd <= 16'h0972;
            973: bcd <= 16'h0973;
            974: bcd <= 16'h0974;
            975: bcd <= 16'h0975;
            976: bcd <= 16'h0976;
            977: bcd <= 16'h0977;
            978: bcd <= 16'h0978;
            979: bcd <= 16'h0979;
            980: bcd <= 16'h0980;
            981: bcd <= 16'h0981;
            982: bcd <= 16'h0982;
            983: bcd <= 16'h0983;
            984: bcd <= 16'h0984;
            985: bcd <= 16'h0985;
            986: bcd <= 16'h0986;
            987: bcd <= 16'h0987;
            988: bcd <= 16'h0988;
            989: bcd <= 16'h0989;
            990: bcd <= 16'h0990;
            991: bcd <= 16'h0991;
            992: bcd <= 16'h0992;
            993: bcd <= 16'h0993;
            994: bcd <= 16'h0994;
            995: bcd <= 16'h0995;
            996: bcd <= 16'h0996;
            997: bcd <= 16'h0997;
            998: bcd <= 16'h0998;
            999: bcd <= 16'h0999;
            1000: bcd <= 16'h1000;
            1001: bcd <= 16'h1001;
            1002: bcd <= 16'h1002;
            1003: bcd <= 16'h1003;
            1004: bcd <= 16'h1004;
            1005: bcd <= 16'h1005;
            1006: bcd <= 16'h1006;
            1007: bcd <= 16'h1007;
            1008: bcd <= 16'h1008;
            1009: bcd <= 16'h1009;
            1010: bcd <= 16'h1010;
            1011: bcd <= 16'h1011;
            1012: bcd <= 16'h1012;
            1013: bcd <= 16'h1013;
            1014: bcd <= 16'h1014;
            1015: bcd <= 16'h1015;
            1016: bcd <= 16'h1016;
            1017: bcd <= 16'h1017;
            1018: bcd <= 16'h1018;
            1019: bcd <= 16'h1019;
            1020: bcd <= 16'h1020;
            1021: bcd <= 16'h1021;
            1022: bcd <= 16'h1022;
            1023: bcd <= 16'h1023;
            1024: bcd <= 16'h1024;
            1025: bcd <= 16'h1025;
            1026: bcd <= 16'h1026;
            1027: bcd <= 16'h1027;
            1028: bcd <= 16'h1028;
            1029: bcd <= 16'h1029;
            1030: bcd <= 16'h1030;
            1031: bcd <= 16'h1031;
            1032: bcd <= 16'h1032;
            1033: bcd <= 16'h1033;
            1034: bcd <= 16'h1034;
            1035: bcd <= 16'h1035;
            1036: bcd <= 16'h1036;
            1037: bcd <= 16'h1037;
            1038: bcd <= 16'h1038;
            1039: bcd <= 16'h1039;
            1040: bcd <= 16'h1040;
            1041: bcd <= 16'h1041;
            1042: bcd <= 16'h1042;
            1043: bcd <= 16'h1043;
            1044: bcd <= 16'h1044;
            1045: bcd <= 16'h1045;
            1046: bcd <= 16'h1046;
            1047: bcd <= 16'h1047;
            1048: bcd <= 16'h1048;
            1049: bcd <= 16'h1049;
            1050: bcd <= 16'h1050;
            1051: bcd <= 16'h1051;
            1052: bcd <= 16'h1052;
            1053: bcd <= 16'h1053;
            1054: bcd <= 16'h1054;
            1055: bcd <= 16'h1055;
            1056: bcd <= 16'h1056;
            1057: bcd <= 16'h1057;
            1058: bcd <= 16'h1058;
            1059: bcd <= 16'h1059;
            1060: bcd <= 16'h1060;
            1061: bcd <= 16'h1061;
            1062: bcd <= 16'h1062;
            1063: bcd <= 16'h1063;
            1064: bcd <= 16'h1064;
            1065: bcd <= 16'h1065;
            1066: bcd <= 16'h1066;
            1067: bcd <= 16'h1067;
            1068: bcd <= 16'h1068;
            1069: bcd <= 16'h1069;
            1070: bcd <= 16'h1070;
            1071: bcd <= 16'h1071;
            1072: bcd <= 16'h1072;
            1073: bcd <= 16'h1073;
            1074: bcd <= 16'h1074;
            1075: bcd <= 16'h1075;
            1076: bcd <= 16'h1076;
            1077: bcd <= 16'h1077;
            1078: bcd <= 16'h1078;
            1079: bcd <= 16'h1079;
            1080: bcd <= 16'h1080;
            1081: bcd <= 16'h1081;
            1082: bcd <= 16'h1082;
            1083: bcd <= 16'h1083;
            1084: bcd <= 16'h1084;
            1085: bcd <= 16'h1085;
            1086: bcd <= 16'h1086;
            1087: bcd <= 16'h1087;
            1088: bcd <= 16'h1088;
            1089: bcd <= 16'h1089;
            1090: bcd <= 16'h1090;
            1091: bcd <= 16'h1091;
            1092: bcd <= 16'h1092;
            1093: bcd <= 16'h1093;
            1094: bcd <= 16'h1094;
            1095: bcd <= 16'h1095;
            1096: bcd <= 16'h1096;
            1097: bcd <= 16'h1097;
            1098: bcd <= 16'h1098;
            1099: bcd <= 16'h1099;
            1100: bcd <= 16'h1100;
            1101: bcd <= 16'h1101;
            1102: bcd <= 16'h1102;
            1103: bcd <= 16'h1103;
            1104: bcd <= 16'h1104;
            1105: bcd <= 16'h1105;
            1106: bcd <= 16'h1106;
            1107: bcd <= 16'h1107;
            1108: bcd <= 16'h1108;
            1109: bcd <= 16'h1109;
            1110: bcd <= 16'h1110;
            1111: bcd <= 16'h1111;
            1112: bcd <= 16'h1112;
            1113: bcd <= 16'h1113;
            1114: bcd <= 16'h1114;
            1115: bcd <= 16'h1115;
            1116: bcd <= 16'h1116;
            1117: bcd <= 16'h1117;
            1118: bcd <= 16'h1118;
            1119: bcd <= 16'h1119;
            1120: bcd <= 16'h1120;
            1121: bcd <= 16'h1121;
            1122: bcd <= 16'h1122;
            1123: bcd <= 16'h1123;
            1124: bcd <= 16'h1124;
            1125: bcd <= 16'h1125;
            1126: bcd <= 16'h1126;
            1127: bcd <= 16'h1127;
            1128: bcd <= 16'h1128;
            1129: bcd <= 16'h1129;
            1130: bcd <= 16'h1130;
            1131: bcd <= 16'h1131;
            1132: bcd <= 16'h1132;
            1133: bcd <= 16'h1133;
            1134: bcd <= 16'h1134;
            1135: bcd <= 16'h1135;
            1136: bcd <= 16'h1136;
            1137: bcd <= 16'h1137;
            1138: bcd <= 16'h1138;
            1139: bcd <= 16'h1139;
            1140: bcd <= 16'h1140;
            1141: bcd <= 16'h1141;
            1142: bcd <= 16'h1142;
            1143: bcd <= 16'h1143;
            1144: bcd <= 16'h1144;
            1145: bcd <= 16'h1145;
            1146: bcd <= 16'h1146;
            1147: bcd <= 16'h1147;
            1148: bcd <= 16'h1148;
            1149: bcd <= 16'h1149;
            1150: bcd <= 16'h1150;
            1151: bcd <= 16'h1151;
            1152: bcd <= 16'h1152;
            1153: bcd <= 16'h1153;
            1154: bcd <= 16'h1154;
            1155: bcd <= 16'h1155;
            1156: bcd <= 16'h1156;
            1157: bcd <= 16'h1157;
            1158: bcd <= 16'h1158;
            1159: bcd <= 16'h1159;
            1160: bcd <= 16'h1160;
            1161: bcd <= 16'h1161;
            1162: bcd <= 16'h1162;
            1163: bcd <= 16'h1163;
            1164: bcd <= 16'h1164;
            1165: bcd <= 16'h1165;
            1166: bcd <= 16'h1166;
            1167: bcd <= 16'h1167;
            1168: bcd <= 16'h1168;
            1169: bcd <= 16'h1169;
            1170: bcd <= 16'h1170;
            1171: bcd <= 16'h1171;
            1172: bcd <= 16'h1172;
            1173: bcd <= 16'h1173;
            1174: bcd <= 16'h1174;
            1175: bcd <= 16'h1175;
            1176: bcd <= 16'h1176;
            1177: bcd <= 16'h1177;
            1178: bcd <= 16'h1178;
            1179: bcd <= 16'h1179;
            1180: bcd <= 16'h1180;
            1181: bcd <= 16'h1181;
            1182: bcd <= 16'h1182;
            1183: bcd <= 16'h1183;
            1184: bcd <= 16'h1184;
            1185: bcd <= 16'h1185;
            1186: bcd <= 16'h1186;
            1187: bcd <= 16'h1187;
            1188: bcd <= 16'h1188;
            1189: bcd <= 16'h1189;
            1190: bcd <= 16'h1190;
            1191: bcd <= 16'h1191;
            1192: bcd <= 16'h1192;
            1193: bcd <= 16'h1193;
            1194: bcd <= 16'h1194;
            1195: bcd <= 16'h1195;
            1196: bcd <= 16'h1196;
            1197: bcd <= 16'h1197;
            1198: bcd <= 16'h1198;
            1199: bcd <= 16'h1199;
            1200: bcd <= 16'h1200;
            1201: bcd <= 16'h1201;
            1202: bcd <= 16'h1202;
            1203: bcd <= 16'h1203;
            1204: bcd <= 16'h1204;
            1205: bcd <= 16'h1205;
            1206: bcd <= 16'h1206;
            1207: bcd <= 16'h1207;
            1208: bcd <= 16'h1208;
            1209: bcd <= 16'h1209;
            1210: bcd <= 16'h1210;
            1211: bcd <= 16'h1211;
            1212: bcd <= 16'h1212;
            1213: bcd <= 16'h1213;
            1214: bcd <= 16'h1214;
            1215: bcd <= 16'h1215;
            1216: bcd <= 16'h1216;
            1217: bcd <= 16'h1217;
            1218: bcd <= 16'h1218;
            1219: bcd <= 16'h1219;
            1220: bcd <= 16'h1220;
            1221: bcd <= 16'h1221;
            1222: bcd <= 16'h1222;
            1223: bcd <= 16'h1223;
            1224: bcd <= 16'h1224;
            1225: bcd <= 16'h1225;
            1226: bcd <= 16'h1226;
            1227: bcd <= 16'h1227;
            1228: bcd <= 16'h1228;
            1229: bcd <= 16'h1229;
            1230: bcd <= 16'h1230;
            1231: bcd <= 16'h1231;
            1232: bcd <= 16'h1232;
            1233: bcd <= 16'h1233;
            1234: bcd <= 16'h1234;
            1235: bcd <= 16'h1235;
            1236: bcd <= 16'h1236;
            1237: bcd <= 16'h1237;
            1238: bcd <= 16'h1238;
            1239: bcd <= 16'h1239;
            1240: bcd <= 16'h1240;
            1241: bcd <= 16'h1241;
            1242: bcd <= 16'h1242;
            1243: bcd <= 16'h1243;
            1244: bcd <= 16'h1244;
            1245: bcd <= 16'h1245;
            1246: bcd <= 16'h1246;
            1247: bcd <= 16'h1247;
            1248: bcd <= 16'h1248;
            1249: bcd <= 16'h1249;
            1250: bcd <= 16'h1250;
            1251: bcd <= 16'h1251;
            1252: bcd <= 16'h1252;
            1253: bcd <= 16'h1253;
            1254: bcd <= 16'h1254;
            1255: bcd <= 16'h1255;
            1256: bcd <= 16'h1256;
            1257: bcd <= 16'h1257;
            1258: bcd <= 16'h1258;
            1259: bcd <= 16'h1259;
            1260: bcd <= 16'h1260;
            1261: bcd <= 16'h1261;
            1262: bcd <= 16'h1262;
            1263: bcd <= 16'h1263;
            1264: bcd <= 16'h1264;
            1265: bcd <= 16'h1265;
            1266: bcd <= 16'h1266;
            1267: bcd <= 16'h1267;
            1268: bcd <= 16'h1268;
            1269: bcd <= 16'h1269;
            1270: bcd <= 16'h1270;
            1271: bcd <= 16'h1271;
            1272: bcd <= 16'h1272;
            1273: bcd <= 16'h1273;
            1274: bcd <= 16'h1274;
            1275: bcd <= 16'h1275;
            1276: bcd <= 16'h1276;
            1277: bcd <= 16'h1277;
            1278: bcd <= 16'h1278;
            1279: bcd <= 16'h1279;
            1280: bcd <= 16'h1280;
            1281: bcd <= 16'h1281;
            1282: bcd <= 16'h1282;
            1283: bcd <= 16'h1283;
            1284: bcd <= 16'h1284;
            1285: bcd <= 16'h1285;
            1286: bcd <= 16'h1286;
            1287: bcd <= 16'h1287;
            1288: bcd <= 16'h1288;
            1289: bcd <= 16'h1289;
            1290: bcd <= 16'h1290;
            1291: bcd <= 16'h1291;
            1292: bcd <= 16'h1292;
            1293: bcd <= 16'h1293;
            1294: bcd <= 16'h1294;
            1295: bcd <= 16'h1295;
            1296: bcd <= 16'h1296;
            1297: bcd <= 16'h1297;
            1298: bcd <= 16'h1298;
            1299: bcd <= 16'h1299;
            1300: bcd <= 16'h1300;
            1301: bcd <= 16'h1301;
            1302: bcd <= 16'h1302;
            1303: bcd <= 16'h1303;
            1304: bcd <= 16'h1304;
            1305: bcd <= 16'h1305;
            1306: bcd <= 16'h1306;
            1307: bcd <= 16'h1307;
            1308: bcd <= 16'h1308;
            1309: bcd <= 16'h1309;
            1310: bcd <= 16'h1310;
            1311: bcd <= 16'h1311;
            1312: bcd <= 16'h1312;
            1313: bcd <= 16'h1313;
            1314: bcd <= 16'h1314;
            1315: bcd <= 16'h1315;
            1316: bcd <= 16'h1316;
            1317: bcd <= 16'h1317;
            1318: bcd <= 16'h1318;
            1319: bcd <= 16'h1319;
            1320: bcd <= 16'h1320;
            1321: bcd <= 16'h1321;
            1322: bcd <= 16'h1322;
            1323: bcd <= 16'h1323;
            1324: bcd <= 16'h1324;
            1325: bcd <= 16'h1325;
            1326: bcd <= 16'h1326;
            1327: bcd <= 16'h1327;
            1328: bcd <= 16'h1328;
            1329: bcd <= 16'h1329;
            1330: bcd <= 16'h1330;
            1331: bcd <= 16'h1331;
            1332: bcd <= 16'h1332;
            1333: bcd <= 16'h1333;
            1334: bcd <= 16'h1334;
            1335: bcd <= 16'h1335;
            1336: bcd <= 16'h1336;
            1337: bcd <= 16'h1337;
            1338: bcd <= 16'h1338;
            1339: bcd <= 16'h1339;
            1340: bcd <= 16'h1340;
            1341: bcd <= 16'h1341;
            1342: bcd <= 16'h1342;
            1343: bcd <= 16'h1343;
            1344: bcd <= 16'h1344;
            1345: bcd <= 16'h1345;
            1346: bcd <= 16'h1346;
            1347: bcd <= 16'h1347;
            1348: bcd <= 16'h1348;
            1349: bcd <= 16'h1349;
            1350: bcd <= 16'h1350;
            1351: bcd <= 16'h1351;
            1352: bcd <= 16'h1352;
            1353: bcd <= 16'h1353;
            1354: bcd <= 16'h1354;
            1355: bcd <= 16'h1355;
            1356: bcd <= 16'h1356;
            1357: bcd <= 16'h1357;
            1358: bcd <= 16'h1358;
            1359: bcd <= 16'h1359;
            1360: bcd <= 16'h1360;
            1361: bcd <= 16'h1361;
            1362: bcd <= 16'h1362;
            1363: bcd <= 16'h1363;
            1364: bcd <= 16'h1364;
            1365: bcd <= 16'h1365;
            1366: bcd <= 16'h1366;
            1367: bcd <= 16'h1367;
            1368: bcd <= 16'h1368;
            1369: bcd <= 16'h1369;
            1370: bcd <= 16'h1370;
            1371: bcd <= 16'h1371;
            1372: bcd <= 16'h1372;
            1373: bcd <= 16'h1373;
            1374: bcd <= 16'h1374;
            1375: bcd <= 16'h1375;
            1376: bcd <= 16'h1376;
            1377: bcd <= 16'h1377;
            1378: bcd <= 16'h1378;
            1379: bcd <= 16'h1379;
            1380: bcd <= 16'h1380;
            1381: bcd <= 16'h1381;
            1382: bcd <= 16'h1382;
            1383: bcd <= 16'h1383;
            1384: bcd <= 16'h1384;
            1385: bcd <= 16'h1385;
            1386: bcd <= 16'h1386;
            1387: bcd <= 16'h1387;
            1388: bcd <= 16'h1388;
            1389: bcd <= 16'h1389;
            1390: bcd <= 16'h1390;
            1391: bcd <= 16'h1391;
            1392: bcd <= 16'h1392;
            1393: bcd <= 16'h1393;
            1394: bcd <= 16'h1394;
            1395: bcd <= 16'h1395;
            1396: bcd <= 16'h1396;
            1397: bcd <= 16'h1397;
            1398: bcd <= 16'h1398;
            1399: bcd <= 16'h1399;
            1400: bcd <= 16'h1400;
            1401: bcd <= 16'h1401;
            1402: bcd <= 16'h1402;
            1403: bcd <= 16'h1403;
            1404: bcd <= 16'h1404;
            1405: bcd <= 16'h1405;
            1406: bcd <= 16'h1406;
            1407: bcd <= 16'h1407;
            1408: bcd <= 16'h1408;
            1409: bcd <= 16'h1409;
            1410: bcd <= 16'h1410;
            1411: bcd <= 16'h1411;
            1412: bcd <= 16'h1412;
            1413: bcd <= 16'h1413;
            1414: bcd <= 16'h1414;
            1415: bcd <= 16'h1415;
            1416: bcd <= 16'h1416;
            1417: bcd <= 16'h1417;
            1418: bcd <= 16'h1418;
            1419: bcd <= 16'h1419;
            1420: bcd <= 16'h1420;
            1421: bcd <= 16'h1421;
            1422: bcd <= 16'h1422;
            1423: bcd <= 16'h1423;
            1424: bcd <= 16'h1424;
            1425: bcd <= 16'h1425;
            1426: bcd <= 16'h1426;
            1427: bcd <= 16'h1427;
            1428: bcd <= 16'h1428;
            1429: bcd <= 16'h1429;
            1430: bcd <= 16'h1430;
            1431: bcd <= 16'h1431;
            1432: bcd <= 16'h1432;
            1433: bcd <= 16'h1433;
            1434: bcd <= 16'h1434;
            1435: bcd <= 16'h1435;
            1436: bcd <= 16'h1436;
            1437: bcd <= 16'h1437;
            1438: bcd <= 16'h1438;
            1439: bcd <= 16'h1439;
            1440: bcd <= 16'h1440;
            1441: bcd <= 16'h1441;
            1442: bcd <= 16'h1442;
            1443: bcd <= 16'h1443;
            1444: bcd <= 16'h1444;
            1445: bcd <= 16'h1445;
            1446: bcd <= 16'h1446;
            1447: bcd <= 16'h1447;
            1448: bcd <= 16'h1448;
            1449: bcd <= 16'h1449;
            1450: bcd <= 16'h1450;
            1451: bcd <= 16'h1451;
            1452: bcd <= 16'h1452;
            1453: bcd <= 16'h1453;
            1454: bcd <= 16'h1454;
            1455: bcd <= 16'h1455;
            1456: bcd <= 16'h1456;
            1457: bcd <= 16'h1457;
            1458: bcd <= 16'h1458;
            1459: bcd <= 16'h1459;
            1460: bcd <= 16'h1460;
            1461: bcd <= 16'h1461;
            1462: bcd <= 16'h1462;
            1463: bcd <= 16'h1463;
            1464: bcd <= 16'h1464;
            1465: bcd <= 16'h1465;
            1466: bcd <= 16'h1466;
            1467: bcd <= 16'h1467;
            1468: bcd <= 16'h1468;
            1469: bcd <= 16'h1469;
            1470: bcd <= 16'h1470;
            1471: bcd <= 16'h1471;
            1472: bcd <= 16'h1472;
            1473: bcd <= 16'h1473;
            1474: bcd <= 16'h1474;
            1475: bcd <= 16'h1475;
            1476: bcd <= 16'h1476;
            1477: bcd <= 16'h1477;
            1478: bcd <= 16'h1478;
            1479: bcd <= 16'h1479;
            1480: bcd <= 16'h1480;
            1481: bcd <= 16'h1481;
            1482: bcd <= 16'h1482;
            1483: bcd <= 16'h1483;
            1484: bcd <= 16'h1484;
            1485: bcd <= 16'h1485;
            1486: bcd <= 16'h1486;
            1487: bcd <= 16'h1487;
            1488: bcd <= 16'h1488;
            1489: bcd <= 16'h1489;
            1490: bcd <= 16'h1490;
            1491: bcd <= 16'h1491;
            1492: bcd <= 16'h1492;
            1493: bcd <= 16'h1493;
            1494: bcd <= 16'h1494;
            1495: bcd <= 16'h1495;
            1496: bcd <= 16'h1496;
            1497: bcd <= 16'h1497;
            1498: bcd <= 16'h1498;
            1499: bcd <= 16'h1499;
            1500: bcd <= 16'h1500;
            1501: bcd <= 16'h1501;
            1502: bcd <= 16'h1502;
            1503: bcd <= 16'h1503;
            1504: bcd <= 16'h1504;
            1505: bcd <= 16'h1505;
            1506: bcd <= 16'h1506;
            1507: bcd <= 16'h1507;
            1508: bcd <= 16'h1508;
            1509: bcd <= 16'h1509;
            1510: bcd <= 16'h1510;
            1511: bcd <= 16'h1511;
            1512: bcd <= 16'h1512;
            1513: bcd <= 16'h1513;
            1514: bcd <= 16'h1514;
            1515: bcd <= 16'h1515;
            1516: bcd <= 16'h1516;
            1517: bcd <= 16'h1517;
            1518: bcd <= 16'h1518;
            1519: bcd <= 16'h1519;
            1520: bcd <= 16'h1520;
            1521: bcd <= 16'h1521;
            1522: bcd <= 16'h1522;
            1523: bcd <= 16'h1523;
            1524: bcd <= 16'h1524;
            1525: bcd <= 16'h1525;
            1526: bcd <= 16'h1526;
            1527: bcd <= 16'h1527;
            1528: bcd <= 16'h1528;
            1529: bcd <= 16'h1529;
            1530: bcd <= 16'h1530;
            1531: bcd <= 16'h1531;
            1532: bcd <= 16'h1532;
            1533: bcd <= 16'h1533;
            1534: bcd <= 16'h1534;
            1535: bcd <= 16'h1535;
            1536: bcd <= 16'h1536;
            1537: bcd <= 16'h1537;
            1538: bcd <= 16'h1538;
            1539: bcd <= 16'h1539;
            1540: bcd <= 16'h1540;
            1541: bcd <= 16'h1541;
            1542: bcd <= 16'h1542;
            1543: bcd <= 16'h1543;
            1544: bcd <= 16'h1544;
            1545: bcd <= 16'h1545;
            1546: bcd <= 16'h1546;
            1547: bcd <= 16'h1547;
            1548: bcd <= 16'h1548;
            1549: bcd <= 16'h1549;
            1550: bcd <= 16'h1550;
            1551: bcd <= 16'h1551;
            1552: bcd <= 16'h1552;
            1553: bcd <= 16'h1553;
            1554: bcd <= 16'h1554;
            1555: bcd <= 16'h1555;
            1556: bcd <= 16'h1556;
            1557: bcd <= 16'h1557;
            1558: bcd <= 16'h1558;
            1559: bcd <= 16'h1559;
            1560: bcd <= 16'h1560;
            1561: bcd <= 16'h1561;
            1562: bcd <= 16'h1562;
            1563: bcd <= 16'h1563;
            1564: bcd <= 16'h1564;
            1565: bcd <= 16'h1565;
            1566: bcd <= 16'h1566;
            1567: bcd <= 16'h1567;
            1568: bcd <= 16'h1568;
            1569: bcd <= 16'h1569;
            1570: bcd <= 16'h1570;
            1571: bcd <= 16'h1571;
            1572: bcd <= 16'h1572;
            1573: bcd <= 16'h1573;
            1574: bcd <= 16'h1574;
            1575: bcd <= 16'h1575;
            1576: bcd <= 16'h1576;
            1577: bcd <= 16'h1577;
            1578: bcd <= 16'h1578;
            1579: bcd <= 16'h1579;
            1580: bcd <= 16'h1580;
            1581: bcd <= 16'h1581;
            1582: bcd <= 16'h1582;
            1583: bcd <= 16'h1583;
            1584: bcd <= 16'h1584;
            1585: bcd <= 16'h1585;
            1586: bcd <= 16'h1586;
            1587: bcd <= 16'h1587;
            1588: bcd <= 16'h1588;
            1589: bcd <= 16'h1589;
            1590: bcd <= 16'h1590;
            1591: bcd <= 16'h1591;
            1592: bcd <= 16'h1592;
            1593: bcd <= 16'h1593;
            1594: bcd <= 16'h1594;
            1595: bcd <= 16'h1595;
            1596: bcd <= 16'h1596;
            1597: bcd <= 16'h1597;
            1598: bcd <= 16'h1598;
            1599: bcd <= 16'h1599;
            1600: bcd <= 16'h1600;
            1601: bcd <= 16'h1601;
            1602: bcd <= 16'h1602;
            1603: bcd <= 16'h1603;
            1604: bcd <= 16'h1604;
            1605: bcd <= 16'h1605;
            1606: bcd <= 16'h1606;
            1607: bcd <= 16'h1607;
            1608: bcd <= 16'h1608;
            1609: bcd <= 16'h1609;
            1610: bcd <= 16'h1610;
            1611: bcd <= 16'h1611;
            1612: bcd <= 16'h1612;
            1613: bcd <= 16'h1613;
            1614: bcd <= 16'h1614;
            1615: bcd <= 16'h1615;
            1616: bcd <= 16'h1616;
            1617: bcd <= 16'h1617;
            1618: bcd <= 16'h1618;
            1619: bcd <= 16'h1619;
            1620: bcd <= 16'h1620;
            1621: bcd <= 16'h1621;
            1622: bcd <= 16'h1622;
            1623: bcd <= 16'h1623;
            1624: bcd <= 16'h1624;
            1625: bcd <= 16'h1625;
            1626: bcd <= 16'h1626;
            1627: bcd <= 16'h1627;
            1628: bcd <= 16'h1628;
            1629: bcd <= 16'h1629;
            1630: bcd <= 16'h1630;
            1631: bcd <= 16'h1631;
            1632: bcd <= 16'h1632;
            1633: bcd <= 16'h1633;
            1634: bcd <= 16'h1634;
            1635: bcd <= 16'h1635;
            1636: bcd <= 16'h1636;
            1637: bcd <= 16'h1637;
            1638: bcd <= 16'h1638;
            1639: bcd <= 16'h1639;
            1640: bcd <= 16'h1640;
            1641: bcd <= 16'h1641;
            1642: bcd <= 16'h1642;
            1643: bcd <= 16'h1643;
            1644: bcd <= 16'h1644;
            1645: bcd <= 16'h1645;
            1646: bcd <= 16'h1646;
            1647: bcd <= 16'h1647;
            1648: bcd <= 16'h1648;
            1649: bcd <= 16'h1649;
            1650: bcd <= 16'h1650;
            1651: bcd <= 16'h1651;
            1652: bcd <= 16'h1652;
            1653: bcd <= 16'h1653;
            1654: bcd <= 16'h1654;
            1655: bcd <= 16'h1655;
            1656: bcd <= 16'h1656;
            1657: bcd <= 16'h1657;
            1658: bcd <= 16'h1658;
            1659: bcd <= 16'h1659;
            1660: bcd <= 16'h1660;
            1661: bcd <= 16'h1661;
            1662: bcd <= 16'h1662;
            1663: bcd <= 16'h1663;
            1664: bcd <= 16'h1664;
            1665: bcd <= 16'h1665;
            1666: bcd <= 16'h1666;
            1667: bcd <= 16'h1667;
            1668: bcd <= 16'h1668;
            1669: bcd <= 16'h1669;
            1670: bcd <= 16'h1670;
            1671: bcd <= 16'h1671;
            1672: bcd <= 16'h1672;
            1673: bcd <= 16'h1673;
            1674: bcd <= 16'h1674;
            1675: bcd <= 16'h1675;
            1676: bcd <= 16'h1676;
            1677: bcd <= 16'h1677;
            1678: bcd <= 16'h1678;
            1679: bcd <= 16'h1679;
            1680: bcd <= 16'h1680;
            1681: bcd <= 16'h1681;
            1682: bcd <= 16'h1682;
            1683: bcd <= 16'h1683;
            1684: bcd <= 16'h1684;
            1685: bcd <= 16'h1685;
            1686: bcd <= 16'h1686;
            1687: bcd <= 16'h1687;
            1688: bcd <= 16'h1688;
            1689: bcd <= 16'h1689;
            1690: bcd <= 16'h1690;
            1691: bcd <= 16'h1691;
            1692: bcd <= 16'h1692;
            1693: bcd <= 16'h1693;
            1694: bcd <= 16'h1694;
            1695: bcd <= 16'h1695;
            1696: bcd <= 16'h1696;
            1697: bcd <= 16'h1697;
            1698: bcd <= 16'h1698;
            1699: bcd <= 16'h1699;
            1700: bcd <= 16'h1700;
            1701: bcd <= 16'h1701;
            1702: bcd <= 16'h1702;
            1703: bcd <= 16'h1703;
            1704: bcd <= 16'h1704;
            1705: bcd <= 16'h1705;
            1706: bcd <= 16'h1706;
            1707: bcd <= 16'h1707;
            1708: bcd <= 16'h1708;
            1709: bcd <= 16'h1709;
            1710: bcd <= 16'h1710;
            1711: bcd <= 16'h1711;
            1712: bcd <= 16'h1712;
            1713: bcd <= 16'h1713;
            1714: bcd <= 16'h1714;
            1715: bcd <= 16'h1715;
            1716: bcd <= 16'h1716;
            1717: bcd <= 16'h1717;
            1718: bcd <= 16'h1718;
            1719: bcd <= 16'h1719;
            1720: bcd <= 16'h1720;
            1721: bcd <= 16'h1721;
            1722: bcd <= 16'h1722;
            1723: bcd <= 16'h1723;
            1724: bcd <= 16'h1724;
            1725: bcd <= 16'h1725;
            1726: bcd <= 16'h1726;
            1727: bcd <= 16'h1727;
            1728: bcd <= 16'h1728;
            1729: bcd <= 16'h1729;
            1730: bcd <= 16'h1730;
            1731: bcd <= 16'h1731;
            1732: bcd <= 16'h1732;
            1733: bcd <= 16'h1733;
            1734: bcd <= 16'h1734;
            1735: bcd <= 16'h1735;
            1736: bcd <= 16'h1736;
            1737: bcd <= 16'h1737;
            1738: bcd <= 16'h1738;
            1739: bcd <= 16'h1739;
            1740: bcd <= 16'h1740;
            1741: bcd <= 16'h1741;
            1742: bcd <= 16'h1742;
            1743: bcd <= 16'h1743;
            1744: bcd <= 16'h1744;
            1745: bcd <= 16'h1745;
            1746: bcd <= 16'h1746;
            1747: bcd <= 16'h1747;
            1748: bcd <= 16'h1748;
            1749: bcd <= 16'h1749;
            1750: bcd <= 16'h1750;
            1751: bcd <= 16'h1751;
            1752: bcd <= 16'h1752;
            1753: bcd <= 16'h1753;
            1754: bcd <= 16'h1754;
            1755: bcd <= 16'h1755;
            1756: bcd <= 16'h1756;
            1757: bcd <= 16'h1757;
            1758: bcd <= 16'h1758;
            1759: bcd <= 16'h1759;
            1760: bcd <= 16'h1760;
            1761: bcd <= 16'h1761;
            1762: bcd <= 16'h1762;
            1763: bcd <= 16'h1763;
            1764: bcd <= 16'h1764;
            1765: bcd <= 16'h1765;
            1766: bcd <= 16'h1766;
            1767: bcd <= 16'h1767;
            1768: bcd <= 16'h1768;
            1769: bcd <= 16'h1769;
            1770: bcd <= 16'h1770;
            1771: bcd <= 16'h1771;
            1772: bcd <= 16'h1772;
            1773: bcd <= 16'h1773;
            1774: bcd <= 16'h1774;
            1775: bcd <= 16'h1775;
            1776: bcd <= 16'h1776;
            1777: bcd <= 16'h1777;
            1778: bcd <= 16'h1778;
            1779: bcd <= 16'h1779;
            1780: bcd <= 16'h1780;
            1781: bcd <= 16'h1781;
            1782: bcd <= 16'h1782;
            1783: bcd <= 16'h1783;
            1784: bcd <= 16'h1784;
            1785: bcd <= 16'h1785;
            1786: bcd <= 16'h1786;
            1787: bcd <= 16'h1787;
            1788: bcd <= 16'h1788;
            1789: bcd <= 16'h1789;
            1790: bcd <= 16'h1790;
            1791: bcd <= 16'h1791;
            1792: bcd <= 16'h1792;
            1793: bcd <= 16'h1793;
            1794: bcd <= 16'h1794;
            1795: bcd <= 16'h1795;
            1796: bcd <= 16'h1796;
            1797: bcd <= 16'h1797;
            1798: bcd <= 16'h1798;
            1799: bcd <= 16'h1799;
            1800: bcd <= 16'h1800;
            1801: bcd <= 16'h1801;
            1802: bcd <= 16'h1802;
            1803: bcd <= 16'h1803;
            1804: bcd <= 16'h1804;
            1805: bcd <= 16'h1805;
            1806: bcd <= 16'h1806;
            1807: bcd <= 16'h1807;
            1808: bcd <= 16'h1808;
            1809: bcd <= 16'h1809;
            1810: bcd <= 16'h1810;
            1811: bcd <= 16'h1811;
            1812: bcd <= 16'h1812;
            1813: bcd <= 16'h1813;
            1814: bcd <= 16'h1814;
            1815: bcd <= 16'h1815;
            1816: bcd <= 16'h1816;
            1817: bcd <= 16'h1817;
            1818: bcd <= 16'h1818;
            1819: bcd <= 16'h1819;
            1820: bcd <= 16'h1820;
            1821: bcd <= 16'h1821;
            1822: bcd <= 16'h1822;
            1823: bcd <= 16'h1823;
            1824: bcd <= 16'h1824;
            1825: bcd <= 16'h1825;
            1826: bcd <= 16'h1826;
            1827: bcd <= 16'h1827;
            1828: bcd <= 16'h1828;
            1829: bcd <= 16'h1829;
            1830: bcd <= 16'h1830;
            1831: bcd <= 16'h1831;
            1832: bcd <= 16'h1832;
            1833: bcd <= 16'h1833;
            1834: bcd <= 16'h1834;
            1835: bcd <= 16'h1835;
            1836: bcd <= 16'h1836;
            1837: bcd <= 16'h1837;
            1838: bcd <= 16'h1838;
            1839: bcd <= 16'h1839;
            1840: bcd <= 16'h1840;
            1841: bcd <= 16'h1841;
            1842: bcd <= 16'h1842;
            1843: bcd <= 16'h1843;
            1844: bcd <= 16'h1844;
            1845: bcd <= 16'h1845;
            1846: bcd <= 16'h1846;
            1847: bcd <= 16'h1847;
            1848: bcd <= 16'h1848;
            1849: bcd <= 16'h1849;
            1850: bcd <= 16'h1850;
            1851: bcd <= 16'h1851;
            1852: bcd <= 16'h1852;
            1853: bcd <= 16'h1853;
            1854: bcd <= 16'h1854;
            1855: bcd <= 16'h1855;
            1856: bcd <= 16'h1856;
            1857: bcd <= 16'h1857;
            1858: bcd <= 16'h1858;
            1859: bcd <= 16'h1859;
            1860: bcd <= 16'h1860;
            1861: bcd <= 16'h1861;
            1862: bcd <= 16'h1862;
            1863: bcd <= 16'h1863;
            1864: bcd <= 16'h1864;
            1865: bcd <= 16'h1865;
            1866: bcd <= 16'h1866;
            1867: bcd <= 16'h1867;
            1868: bcd <= 16'h1868;
            1869: bcd <= 16'h1869;
            1870: bcd <= 16'h1870;
            1871: bcd <= 16'h1871;
            1872: bcd <= 16'h1872;
            1873: bcd <= 16'h1873;
            1874: bcd <= 16'h1874;
            1875: bcd <= 16'h1875;
            1876: bcd <= 16'h1876;
            1877: bcd <= 16'h1877;
            1878: bcd <= 16'h1878;
            1879: bcd <= 16'h1879;
            1880: bcd <= 16'h1880;
            1881: bcd <= 16'h1881;
            1882: bcd <= 16'h1882;
            1883: bcd <= 16'h1883;
            1884: bcd <= 16'h1884;
            1885: bcd <= 16'h1885;
            1886: bcd <= 16'h1886;
            1887: bcd <= 16'h1887;
            1888: bcd <= 16'h1888;
            1889: bcd <= 16'h1889;
            1890: bcd <= 16'h1890;
            1891: bcd <= 16'h1891;
            1892: bcd <= 16'h1892;
            1893: bcd <= 16'h1893;
            1894: bcd <= 16'h1894;
            1895: bcd <= 16'h1895;
            1896: bcd <= 16'h1896;
            1897: bcd <= 16'h1897;
            1898: bcd <= 16'h1898;
            1899: bcd <= 16'h1899;
            1900: bcd <= 16'h1900;
            1901: bcd <= 16'h1901;
            1902: bcd <= 16'h1902;
            1903: bcd <= 16'h1903;
            1904: bcd <= 16'h1904;
            1905: bcd <= 16'h1905;
            1906: bcd <= 16'h1906;
            1907: bcd <= 16'h1907;
            1908: bcd <= 16'h1908;
            1909: bcd <= 16'h1909;
            1910: bcd <= 16'h1910;
            1911: bcd <= 16'h1911;
            1912: bcd <= 16'h1912;
            1913: bcd <= 16'h1913;
            1914: bcd <= 16'h1914;
            1915: bcd <= 16'h1915;
            1916: bcd <= 16'h1916;
            1917: bcd <= 16'h1917;
            1918: bcd <= 16'h1918;
            1919: bcd <= 16'h1919;
            1920: bcd <= 16'h1920;
            1921: bcd <= 16'h1921;
            1922: bcd <= 16'h1922;
            1923: bcd <= 16'h1923;
            1924: bcd <= 16'h1924;
            1925: bcd <= 16'h1925;
            1926: bcd <= 16'h1926;
            1927: bcd <= 16'h1927;
            1928: bcd <= 16'h1928;
            1929: bcd <= 16'h1929;
            1930: bcd <= 16'h1930;
            1931: bcd <= 16'h1931;
            1932: bcd <= 16'h1932;
            1933: bcd <= 16'h1933;
            1934: bcd <= 16'h1934;
            1935: bcd <= 16'h1935;
            1936: bcd <= 16'h1936;
            1937: bcd <= 16'h1937;
            1938: bcd <= 16'h1938;
            1939: bcd <= 16'h1939;
            1940: bcd <= 16'h1940;
            1941: bcd <= 16'h1941;
            1942: bcd <= 16'h1942;
            1943: bcd <= 16'h1943;
            1944: bcd <= 16'h1944;
            1945: bcd <= 16'h1945;
            1946: bcd <= 16'h1946;
            1947: bcd <= 16'h1947;
            1948: bcd <= 16'h1948;
            1949: bcd <= 16'h1949;
            1950: bcd <= 16'h1950;
            1951: bcd <= 16'h1951;
            1952: bcd <= 16'h1952;
            1953: bcd <= 16'h1953;
            1954: bcd <= 16'h1954;
            1955: bcd <= 16'h1955;
            1956: bcd <= 16'h1956;
            1957: bcd <= 16'h1957;
            1958: bcd <= 16'h1958;
            1959: bcd <= 16'h1959;
            1960: bcd <= 16'h1960;
            1961: bcd <= 16'h1961;
            1962: bcd <= 16'h1962;
            1963: bcd <= 16'h1963;
            1964: bcd <= 16'h1964;
            1965: bcd <= 16'h1965;
            1966: bcd <= 16'h1966;
            1967: bcd <= 16'h1967;
            1968: bcd <= 16'h1968;
            1969: bcd <= 16'h1969;
            1970: bcd <= 16'h1970;
            1971: bcd <= 16'h1971;
            1972: bcd <= 16'h1972;
            1973: bcd <= 16'h1973;
            1974: bcd <= 16'h1974;
            1975: bcd <= 16'h1975;
            1976: bcd <= 16'h1976;
            1977: bcd <= 16'h1977;
            1978: bcd <= 16'h1978;
            1979: bcd <= 16'h1979;
            1980: bcd <= 16'h1980;
            1981: bcd <= 16'h1981;
            1982: bcd <= 16'h1982;
            1983: bcd <= 16'h1983;
            1984: bcd <= 16'h1984;
            1985: bcd <= 16'h1985;
            1986: bcd <= 16'h1986;
            1987: bcd <= 16'h1987;
            1988: bcd <= 16'h1988;
            1989: bcd <= 16'h1989;
            1990: bcd <= 16'h1990;
            1991: bcd <= 16'h1991;
            1992: bcd <= 16'h1992;
            1993: bcd <= 16'h1993;
            1994: bcd <= 16'h1994;
            1995: bcd <= 16'h1995;
            1996: bcd <= 16'h1996;
            1997: bcd <= 16'h1997;
            1998: bcd <= 16'h1998;
            1999: bcd <= 16'h1999;
            2000: bcd <= 16'h2000;
            2001: bcd <= 16'h2001;
            2002: bcd <= 16'h2002;
            2003: bcd <= 16'h2003;
            2004: bcd <= 16'h2004;
            2005: bcd <= 16'h2005;
            2006: bcd <= 16'h2006;
            2007: bcd <= 16'h2007;
            2008: bcd <= 16'h2008;
            2009: bcd <= 16'h2009;
            2010: bcd <= 16'h2010;
            2011: bcd <= 16'h2011;
            2012: bcd <= 16'h2012;
            2013: bcd <= 16'h2013;
            2014: bcd <= 16'h2014;
            2015: bcd <= 16'h2015;
            2016: bcd <= 16'h2016;
            2017: bcd <= 16'h2017;
            2018: bcd <= 16'h2018;
            2019: bcd <= 16'h2019;
            2020: bcd <= 16'h2020;
            2021: bcd <= 16'h2021;
            2022: bcd <= 16'h2022;
            2023: bcd <= 16'h2023;
            2024: bcd <= 16'h2024;
            2025: bcd <= 16'h2025;
            2026: bcd <= 16'h2026;
            2027: bcd <= 16'h2027;
            2028: bcd <= 16'h2028;
            2029: bcd <= 16'h2029;
            2030: bcd <= 16'h2030;
            2031: bcd <= 16'h2031;
            2032: bcd <= 16'h2032;
            2033: bcd <= 16'h2033;
            2034: bcd <= 16'h2034;
            2035: bcd <= 16'h2035;
            2036: bcd <= 16'h2036;
            2037: bcd <= 16'h2037;
            2038: bcd <= 16'h2038;
            2039: bcd <= 16'h2039;
            2040: bcd <= 16'h2040;
            2041: bcd <= 16'h2041;
            2042: bcd <= 16'h2042;
            2043: bcd <= 16'h2043;
            2044: bcd <= 16'h2044;
            2045: bcd <= 16'h2045;
            2046: bcd <= 16'h2046;
            2047: bcd <= 16'h2047;
            2048: bcd <= 16'h2048;
            2049: bcd <= 16'h2049;
            2050: bcd <= 16'h2050;
            2051: bcd <= 16'h2051;
            2052: bcd <= 16'h2052;
            2053: bcd <= 16'h2053;
            2054: bcd <= 16'h2054;
            2055: bcd <= 16'h2055;
            2056: bcd <= 16'h2056;
            2057: bcd <= 16'h2057;
            2058: bcd <= 16'h2058;
            2059: bcd <= 16'h2059;
            2060: bcd <= 16'h2060;
            2061: bcd <= 16'h2061;
            2062: bcd <= 16'h2062;
            2063: bcd <= 16'h2063;
            2064: bcd <= 16'h2064;
            2065: bcd <= 16'h2065;
            2066: bcd <= 16'h2066;
            2067: bcd <= 16'h2067;
            2068: bcd <= 16'h2068;
            2069: bcd <= 16'h2069;
            2070: bcd <= 16'h2070;
            2071: bcd <= 16'h2071;
            2072: bcd <= 16'h2072;
            2073: bcd <= 16'h2073;
            2074: bcd <= 16'h2074;
            2075: bcd <= 16'h2075;
            2076: bcd <= 16'h2076;
            2077: bcd <= 16'h2077;
            2078: bcd <= 16'h2078;
            2079: bcd <= 16'h2079;
            2080: bcd <= 16'h2080;
            2081: bcd <= 16'h2081;
            2082: bcd <= 16'h2082;
            2083: bcd <= 16'h2083;
            2084: bcd <= 16'h2084;
            2085: bcd <= 16'h2085;
            2086: bcd <= 16'h2086;
            2087: bcd <= 16'h2087;
            2088: bcd <= 16'h2088;
            2089: bcd <= 16'h2089;
            2090: bcd <= 16'h2090;
            2091: bcd <= 16'h2091;
            2092: bcd <= 16'h2092;
            2093: bcd <= 16'h2093;
            2094: bcd <= 16'h2094;
            2095: bcd <= 16'h2095;
            2096: bcd <= 16'h2096;
            2097: bcd <= 16'h2097;
            2098: bcd <= 16'h2098;
            2099: bcd <= 16'h2099;
            2100: bcd <= 16'h2100;
            2101: bcd <= 16'h2101;
            2102: bcd <= 16'h2102;
            2103: bcd <= 16'h2103;
            2104: bcd <= 16'h2104;
            2105: bcd <= 16'h2105;
            2106: bcd <= 16'h2106;
            2107: bcd <= 16'h2107;
            2108: bcd <= 16'h2108;
            2109: bcd <= 16'h2109;
            2110: bcd <= 16'h2110;
            2111: bcd <= 16'h2111;
            2112: bcd <= 16'h2112;
            2113: bcd <= 16'h2113;
            2114: bcd <= 16'h2114;
            2115: bcd <= 16'h2115;
            2116: bcd <= 16'h2116;
            2117: bcd <= 16'h2117;
            2118: bcd <= 16'h2118;
            2119: bcd <= 16'h2119;
            2120: bcd <= 16'h2120;
            2121: bcd <= 16'h2121;
            2122: bcd <= 16'h2122;
            2123: bcd <= 16'h2123;
            2124: bcd <= 16'h2124;
            2125: bcd <= 16'h2125;
            2126: bcd <= 16'h2126;
            2127: bcd <= 16'h2127;
            2128: bcd <= 16'h2128;
            2129: bcd <= 16'h2129;
            2130: bcd <= 16'h2130;
            2131: bcd <= 16'h2131;
            2132: bcd <= 16'h2132;
            2133: bcd <= 16'h2133;
            2134: bcd <= 16'h2134;
            2135: bcd <= 16'h2135;
            2136: bcd <= 16'h2136;
            2137: bcd <= 16'h2137;
            2138: bcd <= 16'h2138;
            2139: bcd <= 16'h2139;
            2140: bcd <= 16'h2140;
            2141: bcd <= 16'h2141;
            2142: bcd <= 16'h2142;
            2143: bcd <= 16'h2143;
            2144: bcd <= 16'h2144;
            2145: bcd <= 16'h2145;
            2146: bcd <= 16'h2146;
            2147: bcd <= 16'h2147;
            2148: bcd <= 16'h2148;
            2149: bcd <= 16'h2149;
            2150: bcd <= 16'h2150;
            2151: bcd <= 16'h2151;
            2152: bcd <= 16'h2152;
            2153: bcd <= 16'h2153;
            2154: bcd <= 16'h2154;
            2155: bcd <= 16'h2155;
            2156: bcd <= 16'h2156;
            2157: bcd <= 16'h2157;
            2158: bcd <= 16'h2158;
            2159: bcd <= 16'h2159;
            2160: bcd <= 16'h2160;
            2161: bcd <= 16'h2161;
            2162: bcd <= 16'h2162;
            2163: bcd <= 16'h2163;
            2164: bcd <= 16'h2164;
            2165: bcd <= 16'h2165;
            2166: bcd <= 16'h2166;
            2167: bcd <= 16'h2167;
            2168: bcd <= 16'h2168;
            2169: bcd <= 16'h2169;
            2170: bcd <= 16'h2170;
            2171: bcd <= 16'h2171;
            2172: bcd <= 16'h2172;
            2173: bcd <= 16'h2173;
            2174: bcd <= 16'h2174;
            2175: bcd <= 16'h2175;
            2176: bcd <= 16'h2176;
            2177: bcd <= 16'h2177;
            2178: bcd <= 16'h2178;
            2179: bcd <= 16'h2179;
            2180: bcd <= 16'h2180;
            2181: bcd <= 16'h2181;
            2182: bcd <= 16'h2182;
            2183: bcd <= 16'h2183;
            2184: bcd <= 16'h2184;
            2185: bcd <= 16'h2185;
            2186: bcd <= 16'h2186;
            2187: bcd <= 16'h2187;
            2188: bcd <= 16'h2188;
            2189: bcd <= 16'h2189;
            2190: bcd <= 16'h2190;
            2191: bcd <= 16'h2191;
            2192: bcd <= 16'h2192;
            2193: bcd <= 16'h2193;
            2194: bcd <= 16'h2194;
            2195: bcd <= 16'h2195;
            2196: bcd <= 16'h2196;
            2197: bcd <= 16'h2197;
            2198: bcd <= 16'h2198;
            2199: bcd <= 16'h2199;
            2200: bcd <= 16'h2200;
            2201: bcd <= 16'h2201;
            2202: bcd <= 16'h2202;
            2203: bcd <= 16'h2203;
            2204: bcd <= 16'h2204;
            2205: bcd <= 16'h2205;
            2206: bcd <= 16'h2206;
            2207: bcd <= 16'h2207;
            2208: bcd <= 16'h2208;
            2209: bcd <= 16'h2209;
            2210: bcd <= 16'h2210;
            2211: bcd <= 16'h2211;
            2212: bcd <= 16'h2212;
            2213: bcd <= 16'h2213;
            2214: bcd <= 16'h2214;
            2215: bcd <= 16'h2215;
            2216: bcd <= 16'h2216;
            2217: bcd <= 16'h2217;
            2218: bcd <= 16'h2218;
            2219: bcd <= 16'h2219;
            2220: bcd <= 16'h2220;
            2221: bcd <= 16'h2221;
            2222: bcd <= 16'h2222;
            2223: bcd <= 16'h2223;
            2224: bcd <= 16'h2224;
            2225: bcd <= 16'h2225;
            2226: bcd <= 16'h2226;
            2227: bcd <= 16'h2227;
            2228: bcd <= 16'h2228;
            2229: bcd <= 16'h2229;
            2230: bcd <= 16'h2230;
            2231: bcd <= 16'h2231;
            2232: bcd <= 16'h2232;
            2233: bcd <= 16'h2233;
            2234: bcd <= 16'h2234;
            2235: bcd <= 16'h2235;
            2236: bcd <= 16'h2236;
            2237: bcd <= 16'h2237;
            2238: bcd <= 16'h2238;
            2239: bcd <= 16'h2239;
            2240: bcd <= 16'h2240;
            2241: bcd <= 16'h2241;
            2242: bcd <= 16'h2242;
            2243: bcd <= 16'h2243;
            2244: bcd <= 16'h2244;
            2245: bcd <= 16'h2245;
            2246: bcd <= 16'h2246;
            2247: bcd <= 16'h2247;
            2248: bcd <= 16'h2248;
            2249: bcd <= 16'h2249;
            2250: bcd <= 16'h2250;
            2251: bcd <= 16'h2251;
            2252: bcd <= 16'h2252;
            2253: bcd <= 16'h2253;
            2254: bcd <= 16'h2254;
            2255: bcd <= 16'h2255;
            2256: bcd <= 16'h2256;
            2257: bcd <= 16'h2257;
            2258: bcd <= 16'h2258;
            2259: bcd <= 16'h2259;
            2260: bcd <= 16'h2260;
            2261: bcd <= 16'h2261;
            2262: bcd <= 16'h2262;
            2263: bcd <= 16'h2263;
            2264: bcd <= 16'h2264;
            2265: bcd <= 16'h2265;
            2266: bcd <= 16'h2266;
            2267: bcd <= 16'h2267;
            2268: bcd <= 16'h2268;
            2269: bcd <= 16'h2269;
            2270: bcd <= 16'h2270;
            2271: bcd <= 16'h2271;
            2272: bcd <= 16'h2272;
            2273: bcd <= 16'h2273;
            2274: bcd <= 16'h2274;
            2275: bcd <= 16'h2275;
            2276: bcd <= 16'h2276;
            2277: bcd <= 16'h2277;
            2278: bcd <= 16'h2278;
            2279: bcd <= 16'h2279;
            2280: bcd <= 16'h2280;
            2281: bcd <= 16'h2281;
            2282: bcd <= 16'h2282;
            2283: bcd <= 16'h2283;
            2284: bcd <= 16'h2284;
            2285: bcd <= 16'h2285;
            2286: bcd <= 16'h2286;
            2287: bcd <= 16'h2287;
            2288: bcd <= 16'h2288;
            2289: bcd <= 16'h2289;
            2290: bcd <= 16'h2290;
            2291: bcd <= 16'h2291;
            2292: bcd <= 16'h2292;
            2293: bcd <= 16'h2293;
            2294: bcd <= 16'h2294;
            2295: bcd <= 16'h2295;
            2296: bcd <= 16'h2296;
            2297: bcd <= 16'h2297;
            2298: bcd <= 16'h2298;
            2299: bcd <= 16'h2299;
            2300: bcd <= 16'h2300;
            2301: bcd <= 16'h2301;
            2302: bcd <= 16'h2302;
            2303: bcd <= 16'h2303;
            2304: bcd <= 16'h2304;
            2305: bcd <= 16'h2305;
            2306: bcd <= 16'h2306;
            2307: bcd <= 16'h2307;
            2308: bcd <= 16'h2308;
            2309: bcd <= 16'h2309;
            2310: bcd <= 16'h2310;
            2311: bcd <= 16'h2311;
            2312: bcd <= 16'h2312;
            2313: bcd <= 16'h2313;
            2314: bcd <= 16'h2314;
            2315: bcd <= 16'h2315;
            2316: bcd <= 16'h2316;
            2317: bcd <= 16'h2317;
            2318: bcd <= 16'h2318;
            2319: bcd <= 16'h2319;
            2320: bcd <= 16'h2320;
            2321: bcd <= 16'h2321;
            2322: bcd <= 16'h2322;
            2323: bcd <= 16'h2323;
            2324: bcd <= 16'h2324;
            2325: bcd <= 16'h2325;
            2326: bcd <= 16'h2326;
            2327: bcd <= 16'h2327;
            2328: bcd <= 16'h2328;
            2329: bcd <= 16'h2329;
            2330: bcd <= 16'h2330;
            2331: bcd <= 16'h2331;
            2332: bcd <= 16'h2332;
            2333: bcd <= 16'h2333;
            2334: bcd <= 16'h2334;
            2335: bcd <= 16'h2335;
            2336: bcd <= 16'h2336;
            2337: bcd <= 16'h2337;
            2338: bcd <= 16'h2338;
            2339: bcd <= 16'h2339;
            2340: bcd <= 16'h2340;
            2341: bcd <= 16'h2341;
            2342: bcd <= 16'h2342;
            2343: bcd <= 16'h2343;
            2344: bcd <= 16'h2344;
            2345: bcd <= 16'h2345;
            2346: bcd <= 16'h2346;
            2347: bcd <= 16'h2347;
            2348: bcd <= 16'h2348;
            2349: bcd <= 16'h2349;
            2350: bcd <= 16'h2350;
            2351: bcd <= 16'h2351;
            2352: bcd <= 16'h2352;
            2353: bcd <= 16'h2353;
            2354: bcd <= 16'h2354;
            2355: bcd <= 16'h2355;
            2356: bcd <= 16'h2356;
            2357: bcd <= 16'h2357;
            2358: bcd <= 16'h2358;
            2359: bcd <= 16'h2359;
            2360: bcd <= 16'h2360;
            2361: bcd <= 16'h2361;
            2362: bcd <= 16'h2362;
            2363: bcd <= 16'h2363;
            2364: bcd <= 16'h2364;
            2365: bcd <= 16'h2365;
            2366: bcd <= 16'h2366;
            2367: bcd <= 16'h2367;
            2368: bcd <= 16'h2368;
            2369: bcd <= 16'h2369;
            2370: bcd <= 16'h2370;
            2371: bcd <= 16'h2371;
            2372: bcd <= 16'h2372;
            2373: bcd <= 16'h2373;
            2374: bcd <= 16'h2374;
            2375: bcd <= 16'h2375;
            2376: bcd <= 16'h2376;
            2377: bcd <= 16'h2377;
            2378: bcd <= 16'h2378;
            2379: bcd <= 16'h2379;
            2380: bcd <= 16'h2380;
            2381: bcd <= 16'h2381;
            2382: bcd <= 16'h2382;
            2383: bcd <= 16'h2383;
            2384: bcd <= 16'h2384;
            2385: bcd <= 16'h2385;
            2386: bcd <= 16'h2386;
            2387: bcd <= 16'h2387;
            2388: bcd <= 16'h2388;
            2389: bcd <= 16'h2389;
            2390: bcd <= 16'h2390;
            2391: bcd <= 16'h2391;
            2392: bcd <= 16'h2392;
            2393: bcd <= 16'h2393;
            2394: bcd <= 16'h2394;
            2395: bcd <= 16'h2395;
            2396: bcd <= 16'h2396;
            2397: bcd <= 16'h2397;
            2398: bcd <= 16'h2398;
            2399: bcd <= 16'h2399;
            2400: bcd <= 16'h2400;
            2401: bcd <= 16'h2401;
            2402: bcd <= 16'h2402;
            2403: bcd <= 16'h2403;
            2404: bcd <= 16'h2404;
            2405: bcd <= 16'h2405;
            2406: bcd <= 16'h2406;
            2407: bcd <= 16'h2407;
            2408: bcd <= 16'h2408;
            2409: bcd <= 16'h2409;
            2410: bcd <= 16'h2410;
            2411: bcd <= 16'h2411;
            2412: bcd <= 16'h2412;
            2413: bcd <= 16'h2413;
            2414: bcd <= 16'h2414;
            2415: bcd <= 16'h2415;
            2416: bcd <= 16'h2416;
            2417: bcd <= 16'h2417;
            2418: bcd <= 16'h2418;
            2419: bcd <= 16'h2419;
            2420: bcd <= 16'h2420;
            2421: bcd <= 16'h2421;
            2422: bcd <= 16'h2422;
            2423: bcd <= 16'h2423;
            2424: bcd <= 16'h2424;
            2425: bcd <= 16'h2425;
            2426: bcd <= 16'h2426;
            2427: bcd <= 16'h2427;
            2428: bcd <= 16'h2428;
            2429: bcd <= 16'h2429;
            2430: bcd <= 16'h2430;
            2431: bcd <= 16'h2431;
            2432: bcd <= 16'h2432;
            2433: bcd <= 16'h2433;
            2434: bcd <= 16'h2434;
            2435: bcd <= 16'h2435;
            2436: bcd <= 16'h2436;
            2437: bcd <= 16'h2437;
            2438: bcd <= 16'h2438;
            2439: bcd <= 16'h2439;
            2440: bcd <= 16'h2440;
            2441: bcd <= 16'h2441;
            2442: bcd <= 16'h2442;
            2443: bcd <= 16'h2443;
            2444: bcd <= 16'h2444;
            2445: bcd <= 16'h2445;
            2446: bcd <= 16'h2446;
            2447: bcd <= 16'h2447;
            2448: bcd <= 16'h2448;
            2449: bcd <= 16'h2449;
            2450: bcd <= 16'h2450;
            2451: bcd <= 16'h2451;
            2452: bcd <= 16'h2452;
            2453: bcd <= 16'h2453;
            2454: bcd <= 16'h2454;
            2455: bcd <= 16'h2455;
            2456: bcd <= 16'h2456;
            2457: bcd <= 16'h2457;
            2458: bcd <= 16'h2458;
            2459: bcd <= 16'h2459;
            2460: bcd <= 16'h2460;
            2461: bcd <= 16'h2461;
            2462: bcd <= 16'h2462;
            2463: bcd <= 16'h2463;
            2464: bcd <= 16'h2464;
            2465: bcd <= 16'h2465;
            2466: bcd <= 16'h2466;
            2467: bcd <= 16'h2467;
            2468: bcd <= 16'h2468;
            2469: bcd <= 16'h2469;
            2470: bcd <= 16'h2470;
            2471: bcd <= 16'h2471;
            2472: bcd <= 16'h2472;
            2473: bcd <= 16'h2473;
            2474: bcd <= 16'h2474;
            2475: bcd <= 16'h2475;
            2476: bcd <= 16'h2476;
            2477: bcd <= 16'h2477;
            2478: bcd <= 16'h2478;
            2479: bcd <= 16'h2479;
            2480: bcd <= 16'h2480;
            2481: bcd <= 16'h2481;
            2482: bcd <= 16'h2482;
            2483: bcd <= 16'h2483;
            2484: bcd <= 16'h2484;
            2485: bcd <= 16'h2485;
            2486: bcd <= 16'h2486;
            2487: bcd <= 16'h2487;
            2488: bcd <= 16'h2488;
            2489: bcd <= 16'h2489;
            2490: bcd <= 16'h2490;
            2491: bcd <= 16'h2491;
            2492: bcd <= 16'h2492;
            2493: bcd <= 16'h2493;
            2494: bcd <= 16'h2494;
            2495: bcd <= 16'h2495;
            2496: bcd <= 16'h2496;
            2497: bcd <= 16'h2497;
            2498: bcd <= 16'h2498;
            2499: bcd <= 16'h2499;
            2500: bcd <= 16'h2500;
            2501: bcd <= 16'h2501;
            2502: bcd <= 16'h2502;
            2503: bcd <= 16'h2503;
            2504: bcd <= 16'h2504;
            2505: bcd <= 16'h2505;
            2506: bcd <= 16'h2506;
            2507: bcd <= 16'h2507;
            2508: bcd <= 16'h2508;
            2509: bcd <= 16'h2509;
            2510: bcd <= 16'h2510;
            2511: bcd <= 16'h2511;
            2512: bcd <= 16'h2512;
            2513: bcd <= 16'h2513;
            2514: bcd <= 16'h2514;
            2515: bcd <= 16'h2515;
            2516: bcd <= 16'h2516;
            2517: bcd <= 16'h2517;
            2518: bcd <= 16'h2518;
            2519: bcd <= 16'h2519;
            2520: bcd <= 16'h2520;
            2521: bcd <= 16'h2521;
            2522: bcd <= 16'h2522;
            2523: bcd <= 16'h2523;
            2524: bcd <= 16'h2524;
            2525: bcd <= 16'h2525;
            2526: bcd <= 16'h2526;
            2527: bcd <= 16'h2527;
            2528: bcd <= 16'h2528;
            2529: bcd <= 16'h2529;
            2530: bcd <= 16'h2530;
            2531: bcd <= 16'h2531;
            2532: bcd <= 16'h2532;
            2533: bcd <= 16'h2533;
            2534: bcd <= 16'h2534;
            2535: bcd <= 16'h2535;
            2536: bcd <= 16'h2536;
            2537: bcd <= 16'h2537;
            2538: bcd <= 16'h2538;
            2539: bcd <= 16'h2539;
            2540: bcd <= 16'h2540;
            2541: bcd <= 16'h2541;
            2542: bcd <= 16'h2542;
            2543: bcd <= 16'h2543;
            2544: bcd <= 16'h2544;
            2545: bcd <= 16'h2545;
            2546: bcd <= 16'h2546;
            2547: bcd <= 16'h2547;
            2548: bcd <= 16'h2548;
            2549: bcd <= 16'h2549;
            2550: bcd <= 16'h2550;
            2551: bcd <= 16'h2551;
            2552: bcd <= 16'h2552;
            2553: bcd <= 16'h2553;
            2554: bcd <= 16'h2554;
            2555: bcd <= 16'h2555;
            2556: bcd <= 16'h2556;
            2557: bcd <= 16'h2557;
            2558: bcd <= 16'h2558;
            2559: bcd <= 16'h2559;
            2560: bcd <= 16'h2560;
            2561: bcd <= 16'h2561;
            2562: bcd <= 16'h2562;
            2563: bcd <= 16'h2563;
            2564: bcd <= 16'h2564;
            2565: bcd <= 16'h2565;
            2566: bcd <= 16'h2566;
            2567: bcd <= 16'h2567;
            2568: bcd <= 16'h2568;
            2569: bcd <= 16'h2569;
            2570: bcd <= 16'h2570;
            2571: bcd <= 16'h2571;
            2572: bcd <= 16'h2572;
            2573: bcd <= 16'h2573;
            2574: bcd <= 16'h2574;
            2575: bcd <= 16'h2575;
            2576: bcd <= 16'h2576;
            2577: bcd <= 16'h2577;
            2578: bcd <= 16'h2578;
            2579: bcd <= 16'h2579;
            2580: bcd <= 16'h2580;
            2581: bcd <= 16'h2581;
            2582: bcd <= 16'h2582;
            2583: bcd <= 16'h2583;
            2584: bcd <= 16'h2584;
            2585: bcd <= 16'h2585;
            2586: bcd <= 16'h2586;
            2587: bcd <= 16'h2587;
            2588: bcd <= 16'h2588;
            2589: bcd <= 16'h2589;
            2590: bcd <= 16'h2590;
            2591: bcd <= 16'h2591;
            2592: bcd <= 16'h2592;
            2593: bcd <= 16'h2593;
            2594: bcd <= 16'h2594;
            2595: bcd <= 16'h2595;
            2596: bcd <= 16'h2596;
            2597: bcd <= 16'h2597;
            2598: bcd <= 16'h2598;
            2599: bcd <= 16'h2599;
            2600: bcd <= 16'h2600;
            2601: bcd <= 16'h2601;
            2602: bcd <= 16'h2602;
            2603: bcd <= 16'h2603;
            2604: bcd <= 16'h2604;
            2605: bcd <= 16'h2605;
            2606: bcd <= 16'h2606;
            2607: bcd <= 16'h2607;
            2608: bcd <= 16'h2608;
            2609: bcd <= 16'h2609;
            2610: bcd <= 16'h2610;
            2611: bcd <= 16'h2611;
            2612: bcd <= 16'h2612;
            2613: bcd <= 16'h2613;
            2614: bcd <= 16'h2614;
            2615: bcd <= 16'h2615;
            2616: bcd <= 16'h2616;
            2617: bcd <= 16'h2617;
            2618: bcd <= 16'h2618;
            2619: bcd <= 16'h2619;
            2620: bcd <= 16'h2620;
            2621: bcd <= 16'h2621;
            2622: bcd <= 16'h2622;
            2623: bcd <= 16'h2623;
            2624: bcd <= 16'h2624;
            2625: bcd <= 16'h2625;
            2626: bcd <= 16'h2626;
            2627: bcd <= 16'h2627;
            2628: bcd <= 16'h2628;
            2629: bcd <= 16'h2629;
            2630: bcd <= 16'h2630;
            2631: bcd <= 16'h2631;
            2632: bcd <= 16'h2632;
            2633: bcd <= 16'h2633;
            2634: bcd <= 16'h2634;
            2635: bcd <= 16'h2635;
            2636: bcd <= 16'h2636;
            2637: bcd <= 16'h2637;
            2638: bcd <= 16'h2638;
            2639: bcd <= 16'h2639;
            2640: bcd <= 16'h2640;
            2641: bcd <= 16'h2641;
            2642: bcd <= 16'h2642;
            2643: bcd <= 16'h2643;
            2644: bcd <= 16'h2644;
            2645: bcd <= 16'h2645;
            2646: bcd <= 16'h2646;
            2647: bcd <= 16'h2647;
            2648: bcd <= 16'h2648;
            2649: bcd <= 16'h2649;
            2650: bcd <= 16'h2650;
            2651: bcd <= 16'h2651;
            2652: bcd <= 16'h2652;
            2653: bcd <= 16'h2653;
            2654: bcd <= 16'h2654;
            2655: bcd <= 16'h2655;
            2656: bcd <= 16'h2656;
            2657: bcd <= 16'h2657;
            2658: bcd <= 16'h2658;
            2659: bcd <= 16'h2659;
            2660: bcd <= 16'h2660;
            2661: bcd <= 16'h2661;
            2662: bcd <= 16'h2662;
            2663: bcd <= 16'h2663;
            2664: bcd <= 16'h2664;
            2665: bcd <= 16'h2665;
            2666: bcd <= 16'h2666;
            2667: bcd <= 16'h2667;
            2668: bcd <= 16'h2668;
            2669: bcd <= 16'h2669;
            2670: bcd <= 16'h2670;
            2671: bcd <= 16'h2671;
            2672: bcd <= 16'h2672;
            2673: bcd <= 16'h2673;
            2674: bcd <= 16'h2674;
            2675: bcd <= 16'h2675;
            2676: bcd <= 16'h2676;
            2677: bcd <= 16'h2677;
            2678: bcd <= 16'h2678;
            2679: bcd <= 16'h2679;
            2680: bcd <= 16'h2680;
            2681: bcd <= 16'h2681;
            2682: bcd <= 16'h2682;
            2683: bcd <= 16'h2683;
            2684: bcd <= 16'h2684;
            2685: bcd <= 16'h2685;
            2686: bcd <= 16'h2686;
            2687: bcd <= 16'h2687;
            2688: bcd <= 16'h2688;
            2689: bcd <= 16'h2689;
            2690: bcd <= 16'h2690;
            2691: bcd <= 16'h2691;
            2692: bcd <= 16'h2692;
            2693: bcd <= 16'h2693;
            2694: bcd <= 16'h2694;
            2695: bcd <= 16'h2695;
            2696: bcd <= 16'h2696;
            2697: bcd <= 16'h2697;
            2698: bcd <= 16'h2698;
            2699: bcd <= 16'h2699;
            2700: bcd <= 16'h2700;
            2701: bcd <= 16'h2701;
            2702: bcd <= 16'h2702;
            2703: bcd <= 16'h2703;
            2704: bcd <= 16'h2704;
            2705: bcd <= 16'h2705;
            2706: bcd <= 16'h2706;
            2707: bcd <= 16'h2707;
            2708: bcd <= 16'h2708;
            2709: bcd <= 16'h2709;
            2710: bcd <= 16'h2710;
            2711: bcd <= 16'h2711;
            2712: bcd <= 16'h2712;
            2713: bcd <= 16'h2713;
            2714: bcd <= 16'h2714;
            2715: bcd <= 16'h2715;
            2716: bcd <= 16'h2716;
            2717: bcd <= 16'h2717;
            2718: bcd <= 16'h2718;
            2719: bcd <= 16'h2719;
            2720: bcd <= 16'h2720;
            2721: bcd <= 16'h2721;
            2722: bcd <= 16'h2722;
            2723: bcd <= 16'h2723;
            2724: bcd <= 16'h2724;
            2725: bcd <= 16'h2725;
            2726: bcd <= 16'h2726;
            2727: bcd <= 16'h2727;
            2728: bcd <= 16'h2728;
            2729: bcd <= 16'h2729;
            2730: bcd <= 16'h2730;
            2731: bcd <= 16'h2731;
            2732: bcd <= 16'h2732;
            2733: bcd <= 16'h2733;
            2734: bcd <= 16'h2734;
            2735: bcd <= 16'h2735;
            2736: bcd <= 16'h2736;
            2737: bcd <= 16'h2737;
            2738: bcd <= 16'h2738;
            2739: bcd <= 16'h2739;
            2740: bcd <= 16'h2740;
            2741: bcd <= 16'h2741;
            2742: bcd <= 16'h2742;
            2743: bcd <= 16'h2743;
            2744: bcd <= 16'h2744;
            2745: bcd <= 16'h2745;
            2746: bcd <= 16'h2746;
            2747: bcd <= 16'h2747;
            2748: bcd <= 16'h2748;
            2749: bcd <= 16'h2749;
            2750: bcd <= 16'h2750;
            2751: bcd <= 16'h2751;
            2752: bcd <= 16'h2752;
            2753: bcd <= 16'h2753;
            2754: bcd <= 16'h2754;
            2755: bcd <= 16'h2755;
            2756: bcd <= 16'h2756;
            2757: bcd <= 16'h2757;
            2758: bcd <= 16'h2758;
            2759: bcd <= 16'h2759;
            2760: bcd <= 16'h2760;
            2761: bcd <= 16'h2761;
            2762: bcd <= 16'h2762;
            2763: bcd <= 16'h2763;
            2764: bcd <= 16'h2764;
            2765: bcd <= 16'h2765;
            2766: bcd <= 16'h2766;
            2767: bcd <= 16'h2767;
            2768: bcd <= 16'h2768;
            2769: bcd <= 16'h2769;
            2770: bcd <= 16'h2770;
            2771: bcd <= 16'h2771;
            2772: bcd <= 16'h2772;
            2773: bcd <= 16'h2773;
            2774: bcd <= 16'h2774;
            2775: bcd <= 16'h2775;
            2776: bcd <= 16'h2776;
            2777: bcd <= 16'h2777;
            2778: bcd <= 16'h2778;
            2779: bcd <= 16'h2779;
            2780: bcd <= 16'h2780;
            2781: bcd <= 16'h2781;
            2782: bcd <= 16'h2782;
            2783: bcd <= 16'h2783;
            2784: bcd <= 16'h2784;
            2785: bcd <= 16'h2785;
            2786: bcd <= 16'h2786;
            2787: bcd <= 16'h2787;
            2788: bcd <= 16'h2788;
            2789: bcd <= 16'h2789;
            2790: bcd <= 16'h2790;
            2791: bcd <= 16'h2791;
            2792: bcd <= 16'h2792;
            2793: bcd <= 16'h2793;
            2794: bcd <= 16'h2794;
            2795: bcd <= 16'h2795;
            2796: bcd <= 16'h2796;
            2797: bcd <= 16'h2797;
            2798: bcd <= 16'h2798;
            2799: bcd <= 16'h2799;
            2800: bcd <= 16'h2800;
            2801: bcd <= 16'h2801;
            2802: bcd <= 16'h2802;
            2803: bcd <= 16'h2803;
            2804: bcd <= 16'h2804;
            2805: bcd <= 16'h2805;
            2806: bcd <= 16'h2806;
            2807: bcd <= 16'h2807;
            2808: bcd <= 16'h2808;
            2809: bcd <= 16'h2809;
            2810: bcd <= 16'h2810;
            2811: bcd <= 16'h2811;
            2812: bcd <= 16'h2812;
            2813: bcd <= 16'h2813;
            2814: bcd <= 16'h2814;
            2815: bcd <= 16'h2815;
            2816: bcd <= 16'h2816;
            2817: bcd <= 16'h2817;
            2818: bcd <= 16'h2818;
            2819: bcd <= 16'h2819;
            2820: bcd <= 16'h2820;
            2821: bcd <= 16'h2821;
            2822: bcd <= 16'h2822;
            2823: bcd <= 16'h2823;
            2824: bcd <= 16'h2824;
            2825: bcd <= 16'h2825;
            2826: bcd <= 16'h2826;
            2827: bcd <= 16'h2827;
            2828: bcd <= 16'h2828;
            2829: bcd <= 16'h2829;
            2830: bcd <= 16'h2830;
            2831: bcd <= 16'h2831;
            2832: bcd <= 16'h2832;
            2833: bcd <= 16'h2833;
            2834: bcd <= 16'h2834;
            2835: bcd <= 16'h2835;
            2836: bcd <= 16'h2836;
            2837: bcd <= 16'h2837;
            2838: bcd <= 16'h2838;
            2839: bcd <= 16'h2839;
            2840: bcd <= 16'h2840;
            2841: bcd <= 16'h2841;
            2842: bcd <= 16'h2842;
            2843: bcd <= 16'h2843;
            2844: bcd <= 16'h2844;
            2845: bcd <= 16'h2845;
            2846: bcd <= 16'h2846;
            2847: bcd <= 16'h2847;
            2848: bcd <= 16'h2848;
            2849: bcd <= 16'h2849;
            2850: bcd <= 16'h2850;
            2851: bcd <= 16'h2851;
            2852: bcd <= 16'h2852;
            2853: bcd <= 16'h2853;
            2854: bcd <= 16'h2854;
            2855: bcd <= 16'h2855;
            2856: bcd <= 16'h2856;
            2857: bcd <= 16'h2857;
            2858: bcd <= 16'h2858;
            2859: bcd <= 16'h2859;
            2860: bcd <= 16'h2860;
            2861: bcd <= 16'h2861;
            2862: bcd <= 16'h2862;
            2863: bcd <= 16'h2863;
            2864: bcd <= 16'h2864;
            2865: bcd <= 16'h2865;
            2866: bcd <= 16'h2866;
            2867: bcd <= 16'h2867;
            2868: bcd <= 16'h2868;
            2869: bcd <= 16'h2869;
            2870: bcd <= 16'h2870;
            2871: bcd <= 16'h2871;
            2872: bcd <= 16'h2872;
            2873: bcd <= 16'h2873;
            2874: bcd <= 16'h2874;
            2875: bcd <= 16'h2875;
            2876: bcd <= 16'h2876;
            2877: bcd <= 16'h2877;
            2878: bcd <= 16'h2878;
            2879: bcd <= 16'h2879;
            2880: bcd <= 16'h2880;
            2881: bcd <= 16'h2881;
            2882: bcd <= 16'h2882;
            2883: bcd <= 16'h2883;
            2884: bcd <= 16'h2884;
            2885: bcd <= 16'h2885;
            2886: bcd <= 16'h2886;
            2887: bcd <= 16'h2887;
            2888: bcd <= 16'h2888;
            2889: bcd <= 16'h2889;
            2890: bcd <= 16'h2890;
            2891: bcd <= 16'h2891;
            2892: bcd <= 16'h2892;
            2893: bcd <= 16'h2893;
            2894: bcd <= 16'h2894;
            2895: bcd <= 16'h2895;
            2896: bcd <= 16'h2896;
            2897: bcd <= 16'h2897;
            2898: bcd <= 16'h2898;
            2899: bcd <= 16'h2899;
            2900: bcd <= 16'h2900;
            2901: bcd <= 16'h2901;
            2902: bcd <= 16'h2902;
            2903: bcd <= 16'h2903;
            2904: bcd <= 16'h2904;
            2905: bcd <= 16'h2905;
            2906: bcd <= 16'h2906;
            2907: bcd <= 16'h2907;
            2908: bcd <= 16'h2908;
            2909: bcd <= 16'h2909;
            2910: bcd <= 16'h2910;
            2911: bcd <= 16'h2911;
            2912: bcd <= 16'h2912;
            2913: bcd <= 16'h2913;
            2914: bcd <= 16'h2914;
            2915: bcd <= 16'h2915;
            2916: bcd <= 16'h2916;
            2917: bcd <= 16'h2917;
            2918: bcd <= 16'h2918;
            2919: bcd <= 16'h2919;
            2920: bcd <= 16'h2920;
            2921: bcd <= 16'h2921;
            2922: bcd <= 16'h2922;
            2923: bcd <= 16'h2923;
            2924: bcd <= 16'h2924;
            2925: bcd <= 16'h2925;
            2926: bcd <= 16'h2926;
            2927: bcd <= 16'h2927;
            2928: bcd <= 16'h2928;
            2929: bcd <= 16'h2929;
            2930: bcd <= 16'h2930;
            2931: bcd <= 16'h2931;
            2932: bcd <= 16'h2932;
            2933: bcd <= 16'h2933;
            2934: bcd <= 16'h2934;
            2935: bcd <= 16'h2935;
            2936: bcd <= 16'h2936;
            2937: bcd <= 16'h2937;
            2938: bcd <= 16'h2938;
            2939: bcd <= 16'h2939;
            2940: bcd <= 16'h2940;
            2941: bcd <= 16'h2941;
            2942: bcd <= 16'h2942;
            2943: bcd <= 16'h2943;
            2944: bcd <= 16'h2944;
            2945: bcd <= 16'h2945;
            2946: bcd <= 16'h2946;
            2947: bcd <= 16'h2947;
            2948: bcd <= 16'h2948;
            2949: bcd <= 16'h2949;
            2950: bcd <= 16'h2950;
            2951: bcd <= 16'h2951;
            2952: bcd <= 16'h2952;
            2953: bcd <= 16'h2953;
            2954: bcd <= 16'h2954;
            2955: bcd <= 16'h2955;
            2956: bcd <= 16'h2956;
            2957: bcd <= 16'h2957;
            2958: bcd <= 16'h2958;
            2959: bcd <= 16'h2959;
            2960: bcd <= 16'h2960;
            2961: bcd <= 16'h2961;
            2962: bcd <= 16'h2962;
            2963: bcd <= 16'h2963;
            2964: bcd <= 16'h2964;
            2965: bcd <= 16'h2965;
            2966: bcd <= 16'h2966;
            2967: bcd <= 16'h2967;
            2968: bcd <= 16'h2968;
            2969: bcd <= 16'h2969;
            2970: bcd <= 16'h2970;
            2971: bcd <= 16'h2971;
            2972: bcd <= 16'h2972;
            2973: bcd <= 16'h2973;
            2974: bcd <= 16'h2974;
            2975: bcd <= 16'h2975;
            2976: bcd <= 16'h2976;
            2977: bcd <= 16'h2977;
            2978: bcd <= 16'h2978;
            2979: bcd <= 16'h2979;
            2980: bcd <= 16'h2980;
            2981: bcd <= 16'h2981;
            2982: bcd <= 16'h2982;
            2983: bcd <= 16'h2983;
            2984: bcd <= 16'h2984;
            2985: bcd <= 16'h2985;
            2986: bcd <= 16'h2986;
            2987: bcd <= 16'h2987;
            2988: bcd <= 16'h2988;
            2989: bcd <= 16'h2989;
            2990: bcd <= 16'h2990;
            2991: bcd <= 16'h2991;
            2992: bcd <= 16'h2992;
            2993: bcd <= 16'h2993;
            2994: bcd <= 16'h2994;
            2995: bcd <= 16'h2995;
            2996: bcd <= 16'h2996;
            2997: bcd <= 16'h2997;
            2998: bcd <= 16'h2998;
            2999: bcd <= 16'h2999;
            3000: bcd <= 16'h3000;
            3001: bcd <= 16'h3001;
            3002: bcd <= 16'h3002;
            3003: bcd <= 16'h3003;
            3004: bcd <= 16'h3004;
            3005: bcd <= 16'h3005;
            3006: bcd <= 16'h3006;
            3007: bcd <= 16'h3007;
            3008: bcd <= 16'h3008;
            3009: bcd <= 16'h3009;
            3010: bcd <= 16'h3010;
            3011: bcd <= 16'h3011;
            3012: bcd <= 16'h3012;
            3013: bcd <= 16'h3013;
            3014: bcd <= 16'h3014;
            3015: bcd <= 16'h3015;
            3016: bcd <= 16'h3016;
            3017: bcd <= 16'h3017;
            3018: bcd <= 16'h3018;
            3019: bcd <= 16'h3019;
            3020: bcd <= 16'h3020;
            3021: bcd <= 16'h3021;
            3022: bcd <= 16'h3022;
            3023: bcd <= 16'h3023;
            3024: bcd <= 16'h3024;
            3025: bcd <= 16'h3025;
            3026: bcd <= 16'h3026;
            3027: bcd <= 16'h3027;
            3028: bcd <= 16'h3028;
            3029: bcd <= 16'h3029;
            3030: bcd <= 16'h3030;
            3031: bcd <= 16'h3031;
            3032: bcd <= 16'h3032;
            3033: bcd <= 16'h3033;
            3034: bcd <= 16'h3034;
            3035: bcd <= 16'h3035;
            3036: bcd <= 16'h3036;
            3037: bcd <= 16'h3037;
            3038: bcd <= 16'h3038;
            3039: bcd <= 16'h3039;
            3040: bcd <= 16'h3040;
            3041: bcd <= 16'h3041;
            3042: bcd <= 16'h3042;
            3043: bcd <= 16'h3043;
            3044: bcd <= 16'h3044;
            3045: bcd <= 16'h3045;
            3046: bcd <= 16'h3046;
            3047: bcd <= 16'h3047;
            3048: bcd <= 16'h3048;
            3049: bcd <= 16'h3049;
            3050: bcd <= 16'h3050;
            3051: bcd <= 16'h3051;
            3052: bcd <= 16'h3052;
            3053: bcd <= 16'h3053;
            3054: bcd <= 16'h3054;
            3055: bcd <= 16'h3055;
            3056: bcd <= 16'h3056;
            3057: bcd <= 16'h3057;
            3058: bcd <= 16'h3058;
            3059: bcd <= 16'h3059;
            3060: bcd <= 16'h3060;
            3061: bcd <= 16'h3061;
            3062: bcd <= 16'h3062;
            3063: bcd <= 16'h3063;
            3064: bcd <= 16'h3064;
            3065: bcd <= 16'h3065;
            3066: bcd <= 16'h3066;
            3067: bcd <= 16'h3067;
            3068: bcd <= 16'h3068;
            3069: bcd <= 16'h3069;
            3070: bcd <= 16'h3070;
            3071: bcd <= 16'h3071;
            3072: bcd <= 16'h3072;
            3073: bcd <= 16'h3073;
            3074: bcd <= 16'h3074;
            3075: bcd <= 16'h3075;
            3076: bcd <= 16'h3076;
            3077: bcd <= 16'h3077;
            3078: bcd <= 16'h3078;
            3079: bcd <= 16'h3079;
            3080: bcd <= 16'h3080;
            3081: bcd <= 16'h3081;
            3082: bcd <= 16'h3082;
            3083: bcd <= 16'h3083;
            3084: bcd <= 16'h3084;
            3085: bcd <= 16'h3085;
            3086: bcd <= 16'h3086;
            3087: bcd <= 16'h3087;
            3088: bcd <= 16'h3088;
            3089: bcd <= 16'h3089;
            3090: bcd <= 16'h3090;
            3091: bcd <= 16'h3091;
            3092: bcd <= 16'h3092;
            3093: bcd <= 16'h3093;
            3094: bcd <= 16'h3094;
            3095: bcd <= 16'h3095;
            3096: bcd <= 16'h3096;
            3097: bcd <= 16'h3097;
            3098: bcd <= 16'h3098;
            3099: bcd <= 16'h3099;
            3100: bcd <= 16'h3100;
            3101: bcd <= 16'h3101;
            3102: bcd <= 16'h3102;
            3103: bcd <= 16'h3103;
            3104: bcd <= 16'h3104;
            3105: bcd <= 16'h3105;
            3106: bcd <= 16'h3106;
            3107: bcd <= 16'h3107;
            3108: bcd <= 16'h3108;
            3109: bcd <= 16'h3109;
            3110: bcd <= 16'h3110;
            3111: bcd <= 16'h3111;
            3112: bcd <= 16'h3112;
            3113: bcd <= 16'h3113;
            3114: bcd <= 16'h3114;
            3115: bcd <= 16'h3115;
            3116: bcd <= 16'h3116;
            3117: bcd <= 16'h3117;
            3118: bcd <= 16'h3118;
            3119: bcd <= 16'h3119;
            3120: bcd <= 16'h3120;
            3121: bcd <= 16'h3121;
            3122: bcd <= 16'h3122;
            3123: bcd <= 16'h3123;
            3124: bcd <= 16'h3124;
            3125: bcd <= 16'h3125;
            3126: bcd <= 16'h3126;
            3127: bcd <= 16'h3127;
            3128: bcd <= 16'h3128;
            3129: bcd <= 16'h3129;
            3130: bcd <= 16'h3130;
            3131: bcd <= 16'h3131;
            3132: bcd <= 16'h3132;
            3133: bcd <= 16'h3133;
            3134: bcd <= 16'h3134;
            3135: bcd <= 16'h3135;
            3136: bcd <= 16'h3136;
            3137: bcd <= 16'h3137;
            3138: bcd <= 16'h3138;
            3139: bcd <= 16'h3139;
            3140: bcd <= 16'h3140;
            3141: bcd <= 16'h3141;
            3142: bcd <= 16'h3142;
            3143: bcd <= 16'h3143;
            3144: bcd <= 16'h3144;
            3145: bcd <= 16'h3145;
            3146: bcd <= 16'h3146;
            3147: bcd <= 16'h3147;
            3148: bcd <= 16'h3148;
            3149: bcd <= 16'h3149;
            3150: bcd <= 16'h3150;
            3151: bcd <= 16'h3151;
            3152: bcd <= 16'h3152;
            3153: bcd <= 16'h3153;
            3154: bcd <= 16'h3154;
            3155: bcd <= 16'h3155;
            3156: bcd <= 16'h3156;
            3157: bcd <= 16'h3157;
            3158: bcd <= 16'h3158;
            3159: bcd <= 16'h3159;
            3160: bcd <= 16'h3160;
            3161: bcd <= 16'h3161;
            3162: bcd <= 16'h3162;
            3163: bcd <= 16'h3163;
            3164: bcd <= 16'h3164;
            3165: bcd <= 16'h3165;
            3166: bcd <= 16'h3166;
            3167: bcd <= 16'h3167;
            3168: bcd <= 16'h3168;
            3169: bcd <= 16'h3169;
            3170: bcd <= 16'h3170;
            3171: bcd <= 16'h3171;
            3172: bcd <= 16'h3172;
            3173: bcd <= 16'h3173;
            3174: bcd <= 16'h3174;
            3175: bcd <= 16'h3175;
            3176: bcd <= 16'h3176;
            3177: bcd <= 16'h3177;
            3178: bcd <= 16'h3178;
            3179: bcd <= 16'h3179;
            3180: bcd <= 16'h3180;
            3181: bcd <= 16'h3181;
            3182: bcd <= 16'h3182;
            3183: bcd <= 16'h3183;
            3184: bcd <= 16'h3184;
            3185: bcd <= 16'h3185;
            3186: bcd <= 16'h3186;
            3187: bcd <= 16'h3187;
            3188: bcd <= 16'h3188;
            3189: bcd <= 16'h3189;
            3190: bcd <= 16'h3190;
            3191: bcd <= 16'h3191;
            3192: bcd <= 16'h3192;
            3193: bcd <= 16'h3193;
            3194: bcd <= 16'h3194;
            3195: bcd <= 16'h3195;
            3196: bcd <= 16'h3196;
            3197: bcd <= 16'h3197;
            3198: bcd <= 16'h3198;
            3199: bcd <= 16'h3199;
            3200: bcd <= 16'h3200;
            3201: bcd <= 16'h3201;
            3202: bcd <= 16'h3202;
            3203: bcd <= 16'h3203;
            3204: bcd <= 16'h3204;
            3205: bcd <= 16'h3205;
            3206: bcd <= 16'h3206;
            3207: bcd <= 16'h3207;
            3208: bcd <= 16'h3208;
            3209: bcd <= 16'h3209;
            3210: bcd <= 16'h3210;
            3211: bcd <= 16'h3211;
            3212: bcd <= 16'h3212;
            3213: bcd <= 16'h3213;
            3214: bcd <= 16'h3214;
            3215: bcd <= 16'h3215;
            3216: bcd <= 16'h3216;
            3217: bcd <= 16'h3217;
            3218: bcd <= 16'h3218;
            3219: bcd <= 16'h3219;
            3220: bcd <= 16'h3220;
            3221: bcd <= 16'h3221;
            3222: bcd <= 16'h3222;
            3223: bcd <= 16'h3223;
            3224: bcd <= 16'h3224;
            3225: bcd <= 16'h3225;
            3226: bcd <= 16'h3226;
            3227: bcd <= 16'h3227;
            3228: bcd <= 16'h3228;
            3229: bcd <= 16'h3229;
            3230: bcd <= 16'h3230;
            3231: bcd <= 16'h3231;
            3232: bcd <= 16'h3232;
            3233: bcd <= 16'h3233;
            3234: bcd <= 16'h3234;
            3235: bcd <= 16'h3235;
            3236: bcd <= 16'h3236;
            3237: bcd <= 16'h3237;
            3238: bcd <= 16'h3238;
            3239: bcd <= 16'h3239;
            3240: bcd <= 16'h3240;
            3241: bcd <= 16'h3241;
            3242: bcd <= 16'h3242;
            3243: bcd <= 16'h3243;
            3244: bcd <= 16'h3244;
            3245: bcd <= 16'h3245;
            3246: bcd <= 16'h3246;
            3247: bcd <= 16'h3247;
            3248: bcd <= 16'h3248;
            3249: bcd <= 16'h3249;
            3250: bcd <= 16'h3250;
            3251: bcd <= 16'h3251;
            3252: bcd <= 16'h3252;
            3253: bcd <= 16'h3253;
            3254: bcd <= 16'h3254;
            3255: bcd <= 16'h3255;
            3256: bcd <= 16'h3256;
            3257: bcd <= 16'h3257;
            3258: bcd <= 16'h3258;
            3259: bcd <= 16'h3259;
            3260: bcd <= 16'h3260;
            3261: bcd <= 16'h3261;
            3262: bcd <= 16'h3262;
            3263: bcd <= 16'h3263;
            3264: bcd <= 16'h3264;
            3265: bcd <= 16'h3265;
            3266: bcd <= 16'h3266;
            3267: bcd <= 16'h3267;
            3268: bcd <= 16'h3268;
            3269: bcd <= 16'h3269;
            3270: bcd <= 16'h3270;
            3271: bcd <= 16'h3271;
            3272: bcd <= 16'h3272;
            3273: bcd <= 16'h3273;
            3274: bcd <= 16'h3274;
            3275: bcd <= 16'h3275;
            3276: bcd <= 16'h3276;
            3277: bcd <= 16'h3277;
            3278: bcd <= 16'h3278;
            3279: bcd <= 16'h3279;
            3280: bcd <= 16'h3280;
            3281: bcd <= 16'h3281;
            3282: bcd <= 16'h3282;
            3283: bcd <= 16'h3283;
            3284: bcd <= 16'h3284;
            3285: bcd <= 16'h3285;
            3286: bcd <= 16'h3286;
            3287: bcd <= 16'h3287;
            3288: bcd <= 16'h3288;
            3289: bcd <= 16'h3289;
            3290: bcd <= 16'h3290;
            3291: bcd <= 16'h3291;
            3292: bcd <= 16'h3292;
            3293: bcd <= 16'h3293;
            3294: bcd <= 16'h3294;
            3295: bcd <= 16'h3295;
            3296: bcd <= 16'h3296;
            3297: bcd <= 16'h3297;
            3298: bcd <= 16'h3298;
            3299: bcd <= 16'h3299;
            3300: bcd <= 16'h3300;
            3301: bcd <= 16'h3301;
            3302: bcd <= 16'h3302;
            3303: bcd <= 16'h3303;
            3304: bcd <= 16'h3304;
            3305: bcd <= 16'h3305;
            3306: bcd <= 16'h3306;
            3307: bcd <= 16'h3307;
            3308: bcd <= 16'h3308;
            3309: bcd <= 16'h3309;
            3310: bcd <= 16'h3310;
            3311: bcd <= 16'h3311;
            3312: bcd <= 16'h3312;
            3313: bcd <= 16'h3313;
            3314: bcd <= 16'h3314;
            3315: bcd <= 16'h3315;
            3316: bcd <= 16'h3316;
            3317: bcd <= 16'h3317;
            3318: bcd <= 16'h3318;
            3319: bcd <= 16'h3319;
            3320: bcd <= 16'h3320;
            3321: bcd <= 16'h3321;
            3322: bcd <= 16'h3322;
            3323: bcd <= 16'h3323;
            3324: bcd <= 16'h3324;
            3325: bcd <= 16'h3325;
            3326: bcd <= 16'h3326;
            3327: bcd <= 16'h3327;
            3328: bcd <= 16'h3328;
            3329: bcd <= 16'h3329;
            3330: bcd <= 16'h3330;
            3331: bcd <= 16'h3331;
            3332: bcd <= 16'h3332;
            3333: bcd <= 16'h3333;
            3334: bcd <= 16'h3334;
            3335: bcd <= 16'h3335;
            3336: bcd <= 16'h3336;
            3337: bcd <= 16'h3337;
            3338: bcd <= 16'h3338;
            3339: bcd <= 16'h3339;
            3340: bcd <= 16'h3340;
            3341: bcd <= 16'h3341;
            3342: bcd <= 16'h3342;
            3343: bcd <= 16'h3343;
            3344: bcd <= 16'h3344;
            3345: bcd <= 16'h3345;
            3346: bcd <= 16'h3346;
            3347: bcd <= 16'h3347;
            3348: bcd <= 16'h3348;
            3349: bcd <= 16'h3349;
            3350: bcd <= 16'h3350;
            3351: bcd <= 16'h3351;
            3352: bcd <= 16'h3352;
            3353: bcd <= 16'h3353;
            3354: bcd <= 16'h3354;
            3355: bcd <= 16'h3355;
            3356: bcd <= 16'h3356;
            3357: bcd <= 16'h3357;
            3358: bcd <= 16'h3358;
            3359: bcd <= 16'h3359;
            3360: bcd <= 16'h3360;
            3361: bcd <= 16'h3361;
            3362: bcd <= 16'h3362;
            3363: bcd <= 16'h3363;
            3364: bcd <= 16'h3364;
            3365: bcd <= 16'h3365;
            3366: bcd <= 16'h3366;
            3367: bcd <= 16'h3367;
            3368: bcd <= 16'h3368;
            3369: bcd <= 16'h3369;
            3370: bcd <= 16'h3370;
            3371: bcd <= 16'h3371;
            3372: bcd <= 16'h3372;
            3373: bcd <= 16'h3373;
            3374: bcd <= 16'h3374;
            3375: bcd <= 16'h3375;
            3376: bcd <= 16'h3376;
            3377: bcd <= 16'h3377;
            3378: bcd <= 16'h3378;
            3379: bcd <= 16'h3379;
            3380: bcd <= 16'h3380;
            3381: bcd <= 16'h3381;
            3382: bcd <= 16'h3382;
            3383: bcd <= 16'h3383;
            3384: bcd <= 16'h3384;
            3385: bcd <= 16'h3385;
            3386: bcd <= 16'h3386;
            3387: bcd <= 16'h3387;
            3388: bcd <= 16'h3388;
            3389: bcd <= 16'h3389;
            3390: bcd <= 16'h3390;
            3391: bcd <= 16'h3391;
            3392: bcd <= 16'h3392;
            3393: bcd <= 16'h3393;
            3394: bcd <= 16'h3394;
            3395: bcd <= 16'h3395;
            3396: bcd <= 16'h3396;
            3397: bcd <= 16'h3397;
            3398: bcd <= 16'h3398;
            3399: bcd <= 16'h3399;
            3400: bcd <= 16'h3400;
            3401: bcd <= 16'h3401;
            3402: bcd <= 16'h3402;
            3403: bcd <= 16'h3403;
            3404: bcd <= 16'h3404;
            3405: bcd <= 16'h3405;
            3406: bcd <= 16'h3406;
            3407: bcd <= 16'h3407;
            3408: bcd <= 16'h3408;
            3409: bcd <= 16'h3409;
            3410: bcd <= 16'h3410;
            3411: bcd <= 16'h3411;
            3412: bcd <= 16'h3412;
            3413: bcd <= 16'h3413;
            3414: bcd <= 16'h3414;
            3415: bcd <= 16'h3415;
            3416: bcd <= 16'h3416;
            3417: bcd <= 16'h3417;
            3418: bcd <= 16'h3418;
            3419: bcd <= 16'h3419;
            3420: bcd <= 16'h3420;
            3421: bcd <= 16'h3421;
            3422: bcd <= 16'h3422;
            3423: bcd <= 16'h3423;
            3424: bcd <= 16'h3424;
            3425: bcd <= 16'h3425;
            3426: bcd <= 16'h3426;
            3427: bcd <= 16'h3427;
            3428: bcd <= 16'h3428;
            3429: bcd <= 16'h3429;
            3430: bcd <= 16'h3430;
            3431: bcd <= 16'h3431;
            3432: bcd <= 16'h3432;
            3433: bcd <= 16'h3433;
            3434: bcd <= 16'h3434;
            3435: bcd <= 16'h3435;
            3436: bcd <= 16'h3436;
            3437: bcd <= 16'h3437;
            3438: bcd <= 16'h3438;
            3439: bcd <= 16'h3439;
            3440: bcd <= 16'h3440;
            3441: bcd <= 16'h3441;
            3442: bcd <= 16'h3442;
            3443: bcd <= 16'h3443;
            3444: bcd <= 16'h3444;
            3445: bcd <= 16'h3445;
            3446: bcd <= 16'h3446;
            3447: bcd <= 16'h3447;
            3448: bcd <= 16'h3448;
            3449: bcd <= 16'h3449;
            3450: bcd <= 16'h3450;
            3451: bcd <= 16'h3451;
            3452: bcd <= 16'h3452;
            3453: bcd <= 16'h3453;
            3454: bcd <= 16'h3454;
            3455: bcd <= 16'h3455;
            3456: bcd <= 16'h3456;
            3457: bcd <= 16'h3457;
            3458: bcd <= 16'h3458;
            3459: bcd <= 16'h3459;
            3460: bcd <= 16'h3460;
            3461: bcd <= 16'h3461;
            3462: bcd <= 16'h3462;
            3463: bcd <= 16'h3463;
            3464: bcd <= 16'h3464;
            3465: bcd <= 16'h3465;
            3466: bcd <= 16'h3466;
            3467: bcd <= 16'h3467;
            3468: bcd <= 16'h3468;
            3469: bcd <= 16'h3469;
            3470: bcd <= 16'h3470;
            3471: bcd <= 16'h3471;
            3472: bcd <= 16'h3472;
            3473: bcd <= 16'h3473;
            3474: bcd <= 16'h3474;
            3475: bcd <= 16'h3475;
            3476: bcd <= 16'h3476;
            3477: bcd <= 16'h3477;
            3478: bcd <= 16'h3478;
            3479: bcd <= 16'h3479;
            3480: bcd <= 16'h3480;
            3481: bcd <= 16'h3481;
            3482: bcd <= 16'h3482;
            3483: bcd <= 16'h3483;
            3484: bcd <= 16'h3484;
            3485: bcd <= 16'h3485;
            3486: bcd <= 16'h3486;
            3487: bcd <= 16'h3487;
            3488: bcd <= 16'h3488;
            3489: bcd <= 16'h3489;
            3490: bcd <= 16'h3490;
            3491: bcd <= 16'h3491;
            3492: bcd <= 16'h3492;
            3493: bcd <= 16'h3493;
            3494: bcd <= 16'h3494;
            3495: bcd <= 16'h3495;
            3496: bcd <= 16'h3496;
            3497: bcd <= 16'h3497;
            3498: bcd <= 16'h3498;
            3499: bcd <= 16'h3499;
            3500: bcd <= 16'h3500;
            3501: bcd <= 16'h3501;
            3502: bcd <= 16'h3502;
            3503: bcd <= 16'h3503;
            3504: bcd <= 16'h3504;
            3505: bcd <= 16'h3505;
            3506: bcd <= 16'h3506;
            3507: bcd <= 16'h3507;
            3508: bcd <= 16'h3508;
            3509: bcd <= 16'h3509;
            3510: bcd <= 16'h3510;
            3511: bcd <= 16'h3511;
            3512: bcd <= 16'h3512;
            3513: bcd <= 16'h3513;
            3514: bcd <= 16'h3514;
            3515: bcd <= 16'h3515;
            3516: bcd <= 16'h3516;
            3517: bcd <= 16'h3517;
            3518: bcd <= 16'h3518;
            3519: bcd <= 16'h3519;
            3520: bcd <= 16'h3520;
            3521: bcd <= 16'h3521;
            3522: bcd <= 16'h3522;
            3523: bcd <= 16'h3523;
            3524: bcd <= 16'h3524;
            3525: bcd <= 16'h3525;
            3526: bcd <= 16'h3526;
            3527: bcd <= 16'h3527;
            3528: bcd <= 16'h3528;
            3529: bcd <= 16'h3529;
            3530: bcd <= 16'h3530;
            3531: bcd <= 16'h3531;
            3532: bcd <= 16'h3532;
            3533: bcd <= 16'h3533;
            3534: bcd <= 16'h3534;
            3535: bcd <= 16'h3535;
            3536: bcd <= 16'h3536;
            3537: bcd <= 16'h3537;
            3538: bcd <= 16'h3538;
            3539: bcd <= 16'h3539;
            3540: bcd <= 16'h3540;
            3541: bcd <= 16'h3541;
            3542: bcd <= 16'h3542;
            3543: bcd <= 16'h3543;
            3544: bcd <= 16'h3544;
            3545: bcd <= 16'h3545;
            3546: bcd <= 16'h3546;
            3547: bcd <= 16'h3547;
            3548: bcd <= 16'h3548;
            3549: bcd <= 16'h3549;
            3550: bcd <= 16'h3550;
            3551: bcd <= 16'h3551;
            3552: bcd <= 16'h3552;
            3553: bcd <= 16'h3553;
            3554: bcd <= 16'h3554;
            3555: bcd <= 16'h3555;
            3556: bcd <= 16'h3556;
            3557: bcd <= 16'h3557;
            3558: bcd <= 16'h3558;
            3559: bcd <= 16'h3559;
            3560: bcd <= 16'h3560;
            3561: bcd <= 16'h3561;
            3562: bcd <= 16'h3562;
            3563: bcd <= 16'h3563;
            3564: bcd <= 16'h3564;
            3565: bcd <= 16'h3565;
            3566: bcd <= 16'h3566;
            3567: bcd <= 16'h3567;
            3568: bcd <= 16'h3568;
            3569: bcd <= 16'h3569;
            3570: bcd <= 16'h3570;
            3571: bcd <= 16'h3571;
            3572: bcd <= 16'h3572;
            3573: bcd <= 16'h3573;
            3574: bcd <= 16'h3574;
            3575: bcd <= 16'h3575;
            3576: bcd <= 16'h3576;
            3577: bcd <= 16'h3577;
            3578: bcd <= 16'h3578;
            3579: bcd <= 16'h3579;
            3580: bcd <= 16'h3580;
            3581: bcd <= 16'h3581;
            3582: bcd <= 16'h3582;
            3583: bcd <= 16'h3583;
            3584: bcd <= 16'h3584;
            3585: bcd <= 16'h3585;
            3586: bcd <= 16'h3586;
            3587: bcd <= 16'h3587;
            3588: bcd <= 16'h3588;
            3589: bcd <= 16'h3589;
            3590: bcd <= 16'h3590;
            3591: bcd <= 16'h3591;
            3592: bcd <= 16'h3592;
            3593: bcd <= 16'h3593;
            3594: bcd <= 16'h3594;
            3595: bcd <= 16'h3595;
            3596: bcd <= 16'h3596;
            3597: bcd <= 16'h3597;
            3598: bcd <= 16'h3598;
            3599: bcd <= 16'h3599;
            3600: bcd <= 16'h3600;
            3601: bcd <= 16'h3601;
            3602: bcd <= 16'h3602;
            3603: bcd <= 16'h3603;
            3604: bcd <= 16'h3604;
            3605: bcd <= 16'h3605;
            3606: bcd <= 16'h3606;
            3607: bcd <= 16'h3607;
            3608: bcd <= 16'h3608;
            3609: bcd <= 16'h3609;
            3610: bcd <= 16'h3610;
            3611: bcd <= 16'h3611;
            3612: bcd <= 16'h3612;
            3613: bcd <= 16'h3613;
            3614: bcd <= 16'h3614;
            3615: bcd <= 16'h3615;
            3616: bcd <= 16'h3616;
            3617: bcd <= 16'h3617;
            3618: bcd <= 16'h3618;
            3619: bcd <= 16'h3619;
            3620: bcd <= 16'h3620;
            3621: bcd <= 16'h3621;
            3622: bcd <= 16'h3622;
            3623: bcd <= 16'h3623;
            3624: bcd <= 16'h3624;
            3625: bcd <= 16'h3625;
            3626: bcd <= 16'h3626;
            3627: bcd <= 16'h3627;
            3628: bcd <= 16'h3628;
            3629: bcd <= 16'h3629;
            3630: bcd <= 16'h3630;
            3631: bcd <= 16'h3631;
            3632: bcd <= 16'h3632;
            3633: bcd <= 16'h3633;
            3634: bcd <= 16'h3634;
            3635: bcd <= 16'h3635;
            3636: bcd <= 16'h3636;
            3637: bcd <= 16'h3637;
            3638: bcd <= 16'h3638;
            3639: bcd <= 16'h3639;
            3640: bcd <= 16'h3640;
            3641: bcd <= 16'h3641;
            3642: bcd <= 16'h3642;
            3643: bcd <= 16'h3643;
            3644: bcd <= 16'h3644;
            3645: bcd <= 16'h3645;
            3646: bcd <= 16'h3646;
            3647: bcd <= 16'h3647;
            3648: bcd <= 16'h3648;
            3649: bcd <= 16'h3649;
            3650: bcd <= 16'h3650;
            3651: bcd <= 16'h3651;
            3652: bcd <= 16'h3652;
            3653: bcd <= 16'h3653;
            3654: bcd <= 16'h3654;
            3655: bcd <= 16'h3655;
            3656: bcd <= 16'h3656;
            3657: bcd <= 16'h3657;
            3658: bcd <= 16'h3658;
            3659: bcd <= 16'h3659;
            3660: bcd <= 16'h3660;
            3661: bcd <= 16'h3661;
            3662: bcd <= 16'h3662;
            3663: bcd <= 16'h3663;
            3664: bcd <= 16'h3664;
            3665: bcd <= 16'h3665;
            3666: bcd <= 16'h3666;
            3667: bcd <= 16'h3667;
            3668: bcd <= 16'h3668;
            3669: bcd <= 16'h3669;
            3670: bcd <= 16'h3670;
            3671: bcd <= 16'h3671;
            3672: bcd <= 16'h3672;
            3673: bcd <= 16'h3673;
            3674: bcd <= 16'h3674;
            3675: bcd <= 16'h3675;
            3676: bcd <= 16'h3676;
            3677: bcd <= 16'h3677;
            3678: bcd <= 16'h3678;
            3679: bcd <= 16'h3679;
            3680: bcd <= 16'h3680;
            3681: bcd <= 16'h3681;
            3682: bcd <= 16'h3682;
            3683: bcd <= 16'h3683;
            3684: bcd <= 16'h3684;
            3685: bcd <= 16'h3685;
            3686: bcd <= 16'h3686;
            3687: bcd <= 16'h3687;
            3688: bcd <= 16'h3688;
            3689: bcd <= 16'h3689;
            3690: bcd <= 16'h3690;
            3691: bcd <= 16'h3691;
            3692: bcd <= 16'h3692;
            3693: bcd <= 16'h3693;
            3694: bcd <= 16'h3694;
            3695: bcd <= 16'h3695;
            3696: bcd <= 16'h3696;
            3697: bcd <= 16'h3697;
            3698: bcd <= 16'h3698;
            3699: bcd <= 16'h3699;
            3700: bcd <= 16'h3700;
            3701: bcd <= 16'h3701;
            3702: bcd <= 16'h3702;
            3703: bcd <= 16'h3703;
            3704: bcd <= 16'h3704;
            3705: bcd <= 16'h3705;
            3706: bcd <= 16'h3706;
            3707: bcd <= 16'h3707;
            3708: bcd <= 16'h3708;
            3709: bcd <= 16'h3709;
            3710: bcd <= 16'h3710;
            3711: bcd <= 16'h3711;
            3712: bcd <= 16'h3712;
            3713: bcd <= 16'h3713;
            3714: bcd <= 16'h3714;
            3715: bcd <= 16'h3715;
            3716: bcd <= 16'h3716;
            3717: bcd <= 16'h3717;
            3718: bcd <= 16'h3718;
            3719: bcd <= 16'h3719;
            3720: bcd <= 16'h3720;
            3721: bcd <= 16'h3721;
            3722: bcd <= 16'h3722;
            3723: bcd <= 16'h3723;
            3724: bcd <= 16'h3724;
            3725: bcd <= 16'h3725;
            3726: bcd <= 16'h3726;
            3727: bcd <= 16'h3727;
            3728: bcd <= 16'h3728;
            3729: bcd <= 16'h3729;
            3730: bcd <= 16'h3730;
            3731: bcd <= 16'h3731;
            3732: bcd <= 16'h3732;
            3733: bcd <= 16'h3733;
            3734: bcd <= 16'h3734;
            3735: bcd <= 16'h3735;
            3736: bcd <= 16'h3736;
            3737: bcd <= 16'h3737;
            3738: bcd <= 16'h3738;
            3739: bcd <= 16'h3739;
            3740: bcd <= 16'h3740;
            3741: bcd <= 16'h3741;
            3742: bcd <= 16'h3742;
            3743: bcd <= 16'h3743;
            3744: bcd <= 16'h3744;
            3745: bcd <= 16'h3745;
            3746: bcd <= 16'h3746;
            3747: bcd <= 16'h3747;
            3748: bcd <= 16'h3748;
            3749: bcd <= 16'h3749;
            3750: bcd <= 16'h3750;
            3751: bcd <= 16'h3751;
            3752: bcd <= 16'h3752;
            3753: bcd <= 16'h3753;
            3754: bcd <= 16'h3754;
            3755: bcd <= 16'h3755;
            3756: bcd <= 16'h3756;
            3757: bcd <= 16'h3757;
            3758: bcd <= 16'h3758;
            3759: bcd <= 16'h3759;
            3760: bcd <= 16'h3760;
            3761: bcd <= 16'h3761;
            3762: bcd <= 16'h3762;
            3763: bcd <= 16'h3763;
            3764: bcd <= 16'h3764;
            3765: bcd <= 16'h3765;
            3766: bcd <= 16'h3766;
            3767: bcd <= 16'h3767;
            3768: bcd <= 16'h3768;
            3769: bcd <= 16'h3769;
            3770: bcd <= 16'h3770;
            3771: bcd <= 16'h3771;
            3772: bcd <= 16'h3772;
            3773: bcd <= 16'h3773;
            3774: bcd <= 16'h3774;
            3775: bcd <= 16'h3775;
            3776: bcd <= 16'h3776;
            3777: bcd <= 16'h3777;
            3778: bcd <= 16'h3778;
            3779: bcd <= 16'h3779;
            3780: bcd <= 16'h3780;
            3781: bcd <= 16'h3781;
            3782: bcd <= 16'h3782;
            3783: bcd <= 16'h3783;
            3784: bcd <= 16'h3784;
            3785: bcd <= 16'h3785;
            3786: bcd <= 16'h3786;
            3787: bcd <= 16'h3787;
            3788: bcd <= 16'h3788;
            3789: bcd <= 16'h3789;
            3790: bcd <= 16'h3790;
            3791: bcd <= 16'h3791;
            3792: bcd <= 16'h3792;
            3793: bcd <= 16'h3793;
            3794: bcd <= 16'h3794;
            3795: bcd <= 16'h3795;
            3796: bcd <= 16'h3796;
            3797: bcd <= 16'h3797;
            3798: bcd <= 16'h3798;
            3799: bcd <= 16'h3799;
            3800: bcd <= 16'h3800;
            3801: bcd <= 16'h3801;
            3802: bcd <= 16'h3802;
            3803: bcd <= 16'h3803;
            3804: bcd <= 16'h3804;
            3805: bcd <= 16'h3805;
            3806: bcd <= 16'h3806;
            3807: bcd <= 16'h3807;
            3808: bcd <= 16'h3808;
            3809: bcd <= 16'h3809;
            3810: bcd <= 16'h3810;
            3811: bcd <= 16'h3811;
            3812: bcd <= 16'h3812;
            3813: bcd <= 16'h3813;
            3814: bcd <= 16'h3814;
            3815: bcd <= 16'h3815;
            3816: bcd <= 16'h3816;
            3817: bcd <= 16'h3817;
            3818: bcd <= 16'h3818;
            3819: bcd <= 16'h3819;
            3820: bcd <= 16'h3820;
            3821: bcd <= 16'h3821;
            3822: bcd <= 16'h3822;
            3823: bcd <= 16'h3823;
            3824: bcd <= 16'h3824;
            3825: bcd <= 16'h3825;
            3826: bcd <= 16'h3826;
            3827: bcd <= 16'h3827;
            3828: bcd <= 16'h3828;
            3829: bcd <= 16'h3829;
            3830: bcd <= 16'h3830;
            3831: bcd <= 16'h3831;
            3832: bcd <= 16'h3832;
            3833: bcd <= 16'h3833;
            3834: bcd <= 16'h3834;
            3835: bcd <= 16'h3835;
            3836: bcd <= 16'h3836;
            3837: bcd <= 16'h3837;
            3838: bcd <= 16'h3838;
            3839: bcd <= 16'h3839;
            3840: bcd <= 16'h3840;
            3841: bcd <= 16'h3841;
            3842: bcd <= 16'h3842;
            3843: bcd <= 16'h3843;
            3844: bcd <= 16'h3844;
            3845: bcd <= 16'h3845;
            3846: bcd <= 16'h3846;
            3847: bcd <= 16'h3847;
            3848: bcd <= 16'h3848;
            3849: bcd <= 16'h3849;
            3850: bcd <= 16'h3850;
            3851: bcd <= 16'h3851;
            3852: bcd <= 16'h3852;
            3853: bcd <= 16'h3853;
            3854: bcd <= 16'h3854;
            3855: bcd <= 16'h3855;
            3856: bcd <= 16'h3856;
            3857: bcd <= 16'h3857;
            3858: bcd <= 16'h3858;
            3859: bcd <= 16'h3859;
            3860: bcd <= 16'h3860;
            3861: bcd <= 16'h3861;
            3862: bcd <= 16'h3862;
            3863: bcd <= 16'h3863;
            3864: bcd <= 16'h3864;
            3865: bcd <= 16'h3865;
            3866: bcd <= 16'h3866;
            3867: bcd <= 16'h3867;
            3868: bcd <= 16'h3868;
            3869: bcd <= 16'h3869;
            3870: bcd <= 16'h3870;
            3871: bcd <= 16'h3871;
            3872: bcd <= 16'h3872;
            3873: bcd <= 16'h3873;
            3874: bcd <= 16'h3874;
            3875: bcd <= 16'h3875;
            3876: bcd <= 16'h3876;
            3877: bcd <= 16'h3877;
            3878: bcd <= 16'h3878;
            3879: bcd <= 16'h3879;
            3880: bcd <= 16'h3880;
            3881: bcd <= 16'h3881;
            3882: bcd <= 16'h3882;
            3883: bcd <= 16'h3883;
            3884: bcd <= 16'h3884;
            3885: bcd <= 16'h3885;
            3886: bcd <= 16'h3886;
            3887: bcd <= 16'h3887;
            3888: bcd <= 16'h3888;
            3889: bcd <= 16'h3889;
            3890: bcd <= 16'h3890;
            3891: bcd <= 16'h3891;
            3892: bcd <= 16'h3892;
            3893: bcd <= 16'h3893;
            3894: bcd <= 16'h3894;
            3895: bcd <= 16'h3895;
            3896: bcd <= 16'h3896;
            3897: bcd <= 16'h3897;
            3898: bcd <= 16'h3898;
            3899: bcd <= 16'h3899;
            3900: bcd <= 16'h3900;
            3901: bcd <= 16'h3901;
            3902: bcd <= 16'h3902;
            3903: bcd <= 16'h3903;
            3904: bcd <= 16'h3904;
            3905: bcd <= 16'h3905;
            3906: bcd <= 16'h3906;
            3907: bcd <= 16'h3907;
            3908: bcd <= 16'h3908;
            3909: bcd <= 16'h3909;
            3910: bcd <= 16'h3910;
            3911: bcd <= 16'h3911;
            3912: bcd <= 16'h3912;
            3913: bcd <= 16'h3913;
            3914: bcd <= 16'h3914;
            3915: bcd <= 16'h3915;
            3916: bcd <= 16'h3916;
            3917: bcd <= 16'h3917;
            3918: bcd <= 16'h3918;
            3919: bcd <= 16'h3919;
            3920: bcd <= 16'h3920;
            3921: bcd <= 16'h3921;
            3922: bcd <= 16'h3922;
            3923: bcd <= 16'h3923;
            3924: bcd <= 16'h3924;
            3925: bcd <= 16'h3925;
            3926: bcd <= 16'h3926;
            3927: bcd <= 16'h3927;
            3928: bcd <= 16'h3928;
            3929: bcd <= 16'h3929;
            3930: bcd <= 16'h3930;
            3931: bcd <= 16'h3931;
            3932: bcd <= 16'h3932;
            3933: bcd <= 16'h3933;
            3934: bcd <= 16'h3934;
            3935: bcd <= 16'h3935;
            3936: bcd <= 16'h3936;
            3937: bcd <= 16'h3937;
            3938: bcd <= 16'h3938;
            3939: bcd <= 16'h3939;
            3940: bcd <= 16'h3940;
            3941: bcd <= 16'h3941;
            3942: bcd <= 16'h3942;
            3943: bcd <= 16'h3943;
            3944: bcd <= 16'h3944;
            3945: bcd <= 16'h3945;
            3946: bcd <= 16'h3946;
            3947: bcd <= 16'h3947;
            3948: bcd <= 16'h3948;
            3949: bcd <= 16'h3949;
            3950: bcd <= 16'h3950;
            3951: bcd <= 16'h3951;
            3952: bcd <= 16'h3952;
            3953: bcd <= 16'h3953;
            3954: bcd <= 16'h3954;
            3955: bcd <= 16'h3955;
            3956: bcd <= 16'h3956;
            3957: bcd <= 16'h3957;
            3958: bcd <= 16'h3958;
            3959: bcd <= 16'h3959;
            3960: bcd <= 16'h3960;
            3961: bcd <= 16'h3961;
            3962: bcd <= 16'h3962;
            3963: bcd <= 16'h3963;
            3964: bcd <= 16'h3964;
            3965: bcd <= 16'h3965;
            3966: bcd <= 16'h3966;
            3967: bcd <= 16'h3967;
            3968: bcd <= 16'h3968;
            3969: bcd <= 16'h3969;
            3970: bcd <= 16'h3970;
            3971: bcd <= 16'h3971;
            3972: bcd <= 16'h3972;
            3973: bcd <= 16'h3973;
            3974: bcd <= 16'h3974;
            3975: bcd <= 16'h3975;
            3976: bcd <= 16'h3976;
            3977: bcd <= 16'h3977;
            3978: bcd <= 16'h3978;
            3979: bcd <= 16'h3979;
            3980: bcd <= 16'h3980;
            3981: bcd <= 16'h3981;
            3982: bcd <= 16'h3982;
            3983: bcd <= 16'h3983;
            3984: bcd <= 16'h3984;
            3985: bcd <= 16'h3985;
            3986: bcd <= 16'h3986;
            3987: bcd <= 16'h3987;
            3988: bcd <= 16'h3988;
            3989: bcd <= 16'h3989;
            3990: bcd <= 16'h3990;
            3991: bcd <= 16'h3991;
            3992: bcd <= 16'h3992;
            3993: bcd <= 16'h3993;
            3994: bcd <= 16'h3994;
            3995: bcd <= 16'h3995;
            3996: bcd <= 16'h3996;
            3997: bcd <= 16'h3997;
            3998: bcd <= 16'h3998;
            3999: bcd <= 16'h3999;
            4000: bcd <= 16'h4000;
            4001: bcd <= 16'h4001;
            4002: bcd <= 16'h4002;
            4003: bcd <= 16'h4003;
            4004: bcd <= 16'h4004;
            4005: bcd <= 16'h4005;
            4006: bcd <= 16'h4006;
            4007: bcd <= 16'h4007;
            4008: bcd <= 16'h4008;
            4009: bcd <= 16'h4009;
            4010: bcd <= 16'h4010;
            4011: bcd <= 16'h4011;
            4012: bcd <= 16'h4012;
            4013: bcd <= 16'h4013;
            4014: bcd <= 16'h4014;
            4015: bcd <= 16'h4015;
            4016: bcd <= 16'h4016;
            4017: bcd <= 16'h4017;
            4018: bcd <= 16'h4018;
            4019: bcd <= 16'h4019;
            4020: bcd <= 16'h4020;
            4021: bcd <= 16'h4021;
            4022: bcd <= 16'h4022;
            4023: bcd <= 16'h4023;
            4024: bcd <= 16'h4024;
            4025: bcd <= 16'h4025;
            4026: bcd <= 16'h4026;
            4027: bcd <= 16'h4027;
            4028: bcd <= 16'h4028;
            4029: bcd <= 16'h4029;
            4030: bcd <= 16'h4030;
            4031: bcd <= 16'h4031;
            4032: bcd <= 16'h4032;
            4033: bcd <= 16'h4033;
            4034: bcd <= 16'h4034;
            4035: bcd <= 16'h4035;
            4036: bcd <= 16'h4036;
            4037: bcd <= 16'h4037;
            4038: bcd <= 16'h4038;
            4039: bcd <= 16'h4039;
            4040: bcd <= 16'h4040;
            4041: bcd <= 16'h4041;
            4042: bcd <= 16'h4042;
            4043: bcd <= 16'h4043;
            4044: bcd <= 16'h4044;
            4045: bcd <= 16'h4045;
            4046: bcd <= 16'h4046;
            4047: bcd <= 16'h4047;
            4048: bcd <= 16'h4048;
            4049: bcd <= 16'h4049;
            4050: bcd <= 16'h4050;
            4051: bcd <= 16'h4051;
            4052: bcd <= 16'h4052;
            4053: bcd <= 16'h4053;
            4054: bcd <= 16'h4054;
            4055: bcd <= 16'h4055;
            4056: bcd <= 16'h4056;
            4057: bcd <= 16'h4057;
            4058: bcd <= 16'h4058;
            4059: bcd <= 16'h4059;
            4060: bcd <= 16'h4060;
            4061: bcd <= 16'h4061;
            4062: bcd <= 16'h4062;
            4063: bcd <= 16'h4063;
            4064: bcd <= 16'h4064;
            4065: bcd <= 16'h4065;
            4066: bcd <= 16'h4066;
            4067: bcd <= 16'h4067;
            4068: bcd <= 16'h4068;
            4069: bcd <= 16'h4069;
            4070: bcd <= 16'h4070;
            4071: bcd <= 16'h4071;
            4072: bcd <= 16'h4072;
            4073: bcd <= 16'h4073;
            4074: bcd <= 16'h4074;
            4075: bcd <= 16'h4075;
            4076: bcd <= 16'h4076;
            4077: bcd <= 16'h4077;
            4078: bcd <= 16'h4078;
            4079: bcd <= 16'h4079;
            4080: bcd <= 16'h4080;
            4081: bcd <= 16'h4081;
            4082: bcd <= 16'h4082;
            4083: bcd <= 16'h4083;
            4084: bcd <= 16'h4084;
            4085: bcd <= 16'h4085;
            4086: bcd <= 16'h4086;
            4087: bcd <= 16'h4087;
            4088: bcd <= 16'h4088;
            4089: bcd <= 16'h4089;
            4090: bcd <= 16'h4090;
            4091: bcd <= 16'h4091;
            4092: bcd <= 16'h4092;
            4093: bcd <= 16'h4093;
            4094: bcd <= 16'h4094;
            4095: bcd <= 16'h4095;
            4096: bcd <= 16'h4096;
            4097: bcd <= 16'h4097;
            4098: bcd <= 16'h4098;
            4099: bcd <= 16'h4099;
            4100: bcd <= 16'h4100;
            4101: bcd <= 16'h4101;
            4102: bcd <= 16'h4102;
            4103: bcd <= 16'h4103;
            4104: bcd <= 16'h4104;
            4105: bcd <= 16'h4105;
            4106: bcd <= 16'h4106;
            4107: bcd <= 16'h4107;
            4108: bcd <= 16'h4108;
            4109: bcd <= 16'h4109;
            4110: bcd <= 16'h4110;
            4111: bcd <= 16'h4111;
            4112: bcd <= 16'h4112;
            4113: bcd <= 16'h4113;
            4114: bcd <= 16'h4114;
            4115: bcd <= 16'h4115;
            4116: bcd <= 16'h4116;
            4117: bcd <= 16'h4117;
            4118: bcd <= 16'h4118;
            4119: bcd <= 16'h4119;
            4120: bcd <= 16'h4120;
            4121: bcd <= 16'h4121;
            4122: bcd <= 16'h4122;
            4123: bcd <= 16'h4123;
            4124: bcd <= 16'h4124;
            4125: bcd <= 16'h4125;
            4126: bcd <= 16'h4126;
            4127: bcd <= 16'h4127;
            4128: bcd <= 16'h4128;
            4129: bcd <= 16'h4129;
            4130: bcd <= 16'h4130;
            4131: bcd <= 16'h4131;
            4132: bcd <= 16'h4132;
            4133: bcd <= 16'h4133;
            4134: bcd <= 16'h4134;
            4135: bcd <= 16'h4135;
            4136: bcd <= 16'h4136;
            4137: bcd <= 16'h4137;
            4138: bcd <= 16'h4138;
            4139: bcd <= 16'h4139;
            4140: bcd <= 16'h4140;
            4141: bcd <= 16'h4141;
            4142: bcd <= 16'h4142;
            4143: bcd <= 16'h4143;
            4144: bcd <= 16'h4144;
            4145: bcd <= 16'h4145;
            4146: bcd <= 16'h4146;
            4147: bcd <= 16'h4147;
            4148: bcd <= 16'h4148;
            4149: bcd <= 16'h4149;
            4150: bcd <= 16'h4150;
            4151: bcd <= 16'h4151;
            4152: bcd <= 16'h4152;
            4153: bcd <= 16'h4153;
            4154: bcd <= 16'h4154;
            4155: bcd <= 16'h4155;
            4156: bcd <= 16'h4156;
            4157: bcd <= 16'h4157;
            4158: bcd <= 16'h4158;
            4159: bcd <= 16'h4159;
            4160: bcd <= 16'h4160;
            4161: bcd <= 16'h4161;
            4162: bcd <= 16'h4162;
            4163: bcd <= 16'h4163;
            4164: bcd <= 16'h4164;
            4165: bcd <= 16'h4165;
            4166: bcd <= 16'h4166;
            4167: bcd <= 16'h4167;
            4168: bcd <= 16'h4168;
            4169: bcd <= 16'h4169;
            4170: bcd <= 16'h4170;
            4171: bcd <= 16'h4171;
            4172: bcd <= 16'h4172;
            4173: bcd <= 16'h4173;
            4174: bcd <= 16'h4174;
            4175: bcd <= 16'h4175;
            4176: bcd <= 16'h4176;
            4177: bcd <= 16'h4177;
            4178: bcd <= 16'h4178;
            4179: bcd <= 16'h4179;
            4180: bcd <= 16'h4180;
            4181: bcd <= 16'h4181;
            4182: bcd <= 16'h4182;
            4183: bcd <= 16'h4183;
            4184: bcd <= 16'h4184;
            4185: bcd <= 16'h4185;
            4186: bcd <= 16'h4186;
            4187: bcd <= 16'h4187;
            4188: bcd <= 16'h4188;
            4189: bcd <= 16'h4189;
            4190: bcd <= 16'h4190;
            4191: bcd <= 16'h4191;
            4192: bcd <= 16'h4192;
            4193: bcd <= 16'h4193;
            4194: bcd <= 16'h4194;
            4195: bcd <= 16'h4195;
            4196: bcd <= 16'h4196;
            4197: bcd <= 16'h4197;
            4198: bcd <= 16'h4198;
            4199: bcd <= 16'h4199;
            4200: bcd <= 16'h4200;
            4201: bcd <= 16'h4201;
            4202: bcd <= 16'h4202;
            4203: bcd <= 16'h4203;
            4204: bcd <= 16'h4204;
            4205: bcd <= 16'h4205;
            4206: bcd <= 16'h4206;
            4207: bcd <= 16'h4207;
            4208: bcd <= 16'h4208;
            4209: bcd <= 16'h4209;
            4210: bcd <= 16'h4210;
            4211: bcd <= 16'h4211;
            4212: bcd <= 16'h4212;
            4213: bcd <= 16'h4213;
            4214: bcd <= 16'h4214;
            4215: bcd <= 16'h4215;
            4216: bcd <= 16'h4216;
            4217: bcd <= 16'h4217;
            4218: bcd <= 16'h4218;
            4219: bcd <= 16'h4219;
            4220: bcd <= 16'h4220;
            4221: bcd <= 16'h4221;
            4222: bcd <= 16'h4222;
            4223: bcd <= 16'h4223;
            4224: bcd <= 16'h4224;
            4225: bcd <= 16'h4225;
            4226: bcd <= 16'h4226;
            4227: bcd <= 16'h4227;
            4228: bcd <= 16'h4228;
            4229: bcd <= 16'h4229;
            4230: bcd <= 16'h4230;
            4231: bcd <= 16'h4231;
            4232: bcd <= 16'h4232;
            4233: bcd <= 16'h4233;
            4234: bcd <= 16'h4234;
            4235: bcd <= 16'h4235;
            4236: bcd <= 16'h4236;
            4237: bcd <= 16'h4237;
            4238: bcd <= 16'h4238;
            4239: bcd <= 16'h4239;
            4240: bcd <= 16'h4240;
            4241: bcd <= 16'h4241;
            4242: bcd <= 16'h4242;
            4243: bcd <= 16'h4243;
            4244: bcd <= 16'h4244;
            4245: bcd <= 16'h4245;
            4246: bcd <= 16'h4246;
            4247: bcd <= 16'h4247;
            4248: bcd <= 16'h4248;
            4249: bcd <= 16'h4249;
            4250: bcd <= 16'h4250;
            4251: bcd <= 16'h4251;
            4252: bcd <= 16'h4252;
            4253: bcd <= 16'h4253;
            4254: bcd <= 16'h4254;
            4255: bcd <= 16'h4255;
            4256: bcd <= 16'h4256;
            4257: bcd <= 16'h4257;
            4258: bcd <= 16'h4258;
            4259: bcd <= 16'h4259;
            4260: bcd <= 16'h4260;
            4261: bcd <= 16'h4261;
            4262: bcd <= 16'h4262;
            4263: bcd <= 16'h4263;
            4264: bcd <= 16'h4264;
            4265: bcd <= 16'h4265;
            4266: bcd <= 16'h4266;
            4267: bcd <= 16'h4267;
            4268: bcd <= 16'h4268;
            4269: bcd <= 16'h4269;
            4270: bcd <= 16'h4270;
            4271: bcd <= 16'h4271;
            4272: bcd <= 16'h4272;
            4273: bcd <= 16'h4273;
            4274: bcd <= 16'h4274;
            4275: bcd <= 16'h4275;
            4276: bcd <= 16'h4276;
            4277: bcd <= 16'h4277;
            4278: bcd <= 16'h4278;
            4279: bcd <= 16'h4279;
            4280: bcd <= 16'h4280;
            4281: bcd <= 16'h4281;
            4282: bcd <= 16'h4282;
            4283: bcd <= 16'h4283;
            4284: bcd <= 16'h4284;
            4285: bcd <= 16'h4285;
            4286: bcd <= 16'h4286;
            4287: bcd <= 16'h4287;
            4288: bcd <= 16'h4288;
            4289: bcd <= 16'h4289;
            4290: bcd <= 16'h4290;
            4291: bcd <= 16'h4291;
            4292: bcd <= 16'h4292;
            4293: bcd <= 16'h4293;
            4294: bcd <= 16'h4294;
            4295: bcd <= 16'h4295;
            4296: bcd <= 16'h4296;
            4297: bcd <= 16'h4297;
            4298: bcd <= 16'h4298;
            4299: bcd <= 16'h4299;
            4300: bcd <= 16'h4300;
            4301: bcd <= 16'h4301;
            4302: bcd <= 16'h4302;
            4303: bcd <= 16'h4303;
            4304: bcd <= 16'h4304;
            4305: bcd <= 16'h4305;
            4306: bcd <= 16'h4306;
            4307: bcd <= 16'h4307;
            4308: bcd <= 16'h4308;
            4309: bcd <= 16'h4309;
            4310: bcd <= 16'h4310;
            4311: bcd <= 16'h4311;
            4312: bcd <= 16'h4312;
            4313: bcd <= 16'h4313;
            4314: bcd <= 16'h4314;
            4315: bcd <= 16'h4315;
            4316: bcd <= 16'h4316;
            4317: bcd <= 16'h4317;
            4318: bcd <= 16'h4318;
            4319: bcd <= 16'h4319;
            4320: bcd <= 16'h4320;
            4321: bcd <= 16'h4321;
            4322: bcd <= 16'h4322;
            4323: bcd <= 16'h4323;
            4324: bcd <= 16'h4324;
            4325: bcd <= 16'h4325;
            4326: bcd <= 16'h4326;
            4327: bcd <= 16'h4327;
            4328: bcd <= 16'h4328;
            4329: bcd <= 16'h4329;
            4330: bcd <= 16'h4330;
            4331: bcd <= 16'h4331;
            4332: bcd <= 16'h4332;
            4333: bcd <= 16'h4333;
            4334: bcd <= 16'h4334;
            4335: bcd <= 16'h4335;
            4336: bcd <= 16'h4336;
            4337: bcd <= 16'h4337;
            4338: bcd <= 16'h4338;
            4339: bcd <= 16'h4339;
            4340: bcd <= 16'h4340;
            4341: bcd <= 16'h4341;
            4342: bcd <= 16'h4342;
            4343: bcd <= 16'h4343;
            4344: bcd <= 16'h4344;
            4345: bcd <= 16'h4345;
            4346: bcd <= 16'h4346;
            4347: bcd <= 16'h4347;
            4348: bcd <= 16'h4348;
            4349: bcd <= 16'h4349;
            4350: bcd <= 16'h4350;
            4351: bcd <= 16'h4351;
            4352: bcd <= 16'h4352;
            4353: bcd <= 16'h4353;
            4354: bcd <= 16'h4354;
            4355: bcd <= 16'h4355;
            4356: bcd <= 16'h4356;
            4357: bcd <= 16'h4357;
            4358: bcd <= 16'h4358;
            4359: bcd <= 16'h4359;
            4360: bcd <= 16'h4360;
            4361: bcd <= 16'h4361;
            4362: bcd <= 16'h4362;
            4363: bcd <= 16'h4363;
            4364: bcd <= 16'h4364;
            4365: bcd <= 16'h4365;
            4366: bcd <= 16'h4366;
            4367: bcd <= 16'h4367;
            4368: bcd <= 16'h4368;
            4369: bcd <= 16'h4369;
            4370: bcd <= 16'h4370;
            4371: bcd <= 16'h4371;
            4372: bcd <= 16'h4372;
            4373: bcd <= 16'h4373;
            4374: bcd <= 16'h4374;
            4375: bcd <= 16'h4375;
            4376: bcd <= 16'h4376;
            4377: bcd <= 16'h4377;
            4378: bcd <= 16'h4378;
            4379: bcd <= 16'h4379;
            4380: bcd <= 16'h4380;
            4381: bcd <= 16'h4381;
            4382: bcd <= 16'h4382;
            4383: bcd <= 16'h4383;
            4384: bcd <= 16'h4384;
            4385: bcd <= 16'h4385;
            4386: bcd <= 16'h4386;
            4387: bcd <= 16'h4387;
            4388: bcd <= 16'h4388;
            4389: bcd <= 16'h4389;
            4390: bcd <= 16'h4390;
            4391: bcd <= 16'h4391;
            4392: bcd <= 16'h4392;
            4393: bcd <= 16'h4393;
            4394: bcd <= 16'h4394;
            4395: bcd <= 16'h4395;
            4396: bcd <= 16'h4396;
            4397: bcd <= 16'h4397;
            4398: bcd <= 16'h4398;
            4399: bcd <= 16'h4399;
            4400: bcd <= 16'h4400;
            4401: bcd <= 16'h4401;
            4402: bcd <= 16'h4402;
            4403: bcd <= 16'h4403;
            4404: bcd <= 16'h4404;
            4405: bcd <= 16'h4405;
            4406: bcd <= 16'h4406;
            4407: bcd <= 16'h4407;
            4408: bcd <= 16'h4408;
            4409: bcd <= 16'h4409;
            4410: bcd <= 16'h4410;
            4411: bcd <= 16'h4411;
            4412: bcd <= 16'h4412;
            4413: bcd <= 16'h4413;
            4414: bcd <= 16'h4414;
            4415: bcd <= 16'h4415;
            4416: bcd <= 16'h4416;
            4417: bcd <= 16'h4417;
            4418: bcd <= 16'h4418;
            4419: bcd <= 16'h4419;
            4420: bcd <= 16'h4420;
            4421: bcd <= 16'h4421;
            4422: bcd <= 16'h4422;
            4423: bcd <= 16'h4423;
            4424: bcd <= 16'h4424;
            4425: bcd <= 16'h4425;
            4426: bcd <= 16'h4426;
            4427: bcd <= 16'h4427;
            4428: bcd <= 16'h4428;
            4429: bcd <= 16'h4429;
            4430: bcd <= 16'h4430;
            4431: bcd <= 16'h4431;
            4432: bcd <= 16'h4432;
            4433: bcd <= 16'h4433;
            4434: bcd <= 16'h4434;
            4435: bcd <= 16'h4435;
            4436: bcd <= 16'h4436;
            4437: bcd <= 16'h4437;
            4438: bcd <= 16'h4438;
            4439: bcd <= 16'h4439;
            4440: bcd <= 16'h4440;
            4441: bcd <= 16'h4441;
            4442: bcd <= 16'h4442;
            4443: bcd <= 16'h4443;
            4444: bcd <= 16'h4444;
            4445: bcd <= 16'h4445;
            4446: bcd <= 16'h4446;
            4447: bcd <= 16'h4447;
            4448: bcd <= 16'h4448;
            4449: bcd <= 16'h4449;
            4450: bcd <= 16'h4450;
            4451: bcd <= 16'h4451;
            4452: bcd <= 16'h4452;
            4453: bcd <= 16'h4453;
            4454: bcd <= 16'h4454;
            4455: bcd <= 16'h4455;
            4456: bcd <= 16'h4456;
            4457: bcd <= 16'h4457;
            4458: bcd <= 16'h4458;
            4459: bcd <= 16'h4459;
            4460: bcd <= 16'h4460;
            4461: bcd <= 16'h4461;
            4462: bcd <= 16'h4462;
            4463: bcd <= 16'h4463;
            4464: bcd <= 16'h4464;
            4465: bcd <= 16'h4465;
            4466: bcd <= 16'h4466;
            4467: bcd <= 16'h4467;
            4468: bcd <= 16'h4468;
            4469: bcd <= 16'h4469;
            4470: bcd <= 16'h4470;
            4471: bcd <= 16'h4471;
            4472: bcd <= 16'h4472;
            4473: bcd <= 16'h4473;
            4474: bcd <= 16'h4474;
            4475: bcd <= 16'h4475;
            4476: bcd <= 16'h4476;
            4477: bcd <= 16'h4477;
            4478: bcd <= 16'h4478;
            4479: bcd <= 16'h4479;
            4480: bcd <= 16'h4480;
            4481: bcd <= 16'h4481;
            4482: bcd <= 16'h4482;
            4483: bcd <= 16'h4483;
            4484: bcd <= 16'h4484;
            4485: bcd <= 16'h4485;
            4486: bcd <= 16'h4486;
            4487: bcd <= 16'h4487;
            4488: bcd <= 16'h4488;
            4489: bcd <= 16'h4489;
            4490: bcd <= 16'h4490;
            4491: bcd <= 16'h4491;
            4492: bcd <= 16'h4492;
            4493: bcd <= 16'h4493;
            4494: bcd <= 16'h4494;
            4495: bcd <= 16'h4495;
            4496: bcd <= 16'h4496;
            4497: bcd <= 16'h4497;
            4498: bcd <= 16'h4498;
            4499: bcd <= 16'h4499;
            4500: bcd <= 16'h4500;
            4501: bcd <= 16'h4501;
            4502: bcd <= 16'h4502;
            4503: bcd <= 16'h4503;
            4504: bcd <= 16'h4504;
            4505: bcd <= 16'h4505;
            4506: bcd <= 16'h4506;
            4507: bcd <= 16'h4507;
            4508: bcd <= 16'h4508;
            4509: bcd <= 16'h4509;
            4510: bcd <= 16'h4510;
            4511: bcd <= 16'h4511;
            4512: bcd <= 16'h4512;
            4513: bcd <= 16'h4513;
            4514: bcd <= 16'h4514;
            4515: bcd <= 16'h4515;
            4516: bcd <= 16'h4516;
            4517: bcd <= 16'h4517;
            4518: bcd <= 16'h4518;
            4519: bcd <= 16'h4519;
            4520: bcd <= 16'h4520;
            4521: bcd <= 16'h4521;
            4522: bcd <= 16'h4522;
            4523: bcd <= 16'h4523;
            4524: bcd <= 16'h4524;
            4525: bcd <= 16'h4525;
            4526: bcd <= 16'h4526;
            4527: bcd <= 16'h4527;
            4528: bcd <= 16'h4528;
            4529: bcd <= 16'h4529;
            4530: bcd <= 16'h4530;
            4531: bcd <= 16'h4531;
            4532: bcd <= 16'h4532;
            4533: bcd <= 16'h4533;
            4534: bcd <= 16'h4534;
            4535: bcd <= 16'h4535;
            4536: bcd <= 16'h4536;
            4537: bcd <= 16'h4537;
            4538: bcd <= 16'h4538;
            4539: bcd <= 16'h4539;
            4540: bcd <= 16'h4540;
            4541: bcd <= 16'h4541;
            4542: bcd <= 16'h4542;
            4543: bcd <= 16'h4543;
            4544: bcd <= 16'h4544;
            4545: bcd <= 16'h4545;
            4546: bcd <= 16'h4546;
            4547: bcd <= 16'h4547;
            4548: bcd <= 16'h4548;
            4549: bcd <= 16'h4549;
            4550: bcd <= 16'h4550;
            4551: bcd <= 16'h4551;
            4552: bcd <= 16'h4552;
            4553: bcd <= 16'h4553;
            4554: bcd <= 16'h4554;
            4555: bcd <= 16'h4555;
            4556: bcd <= 16'h4556;
            4557: bcd <= 16'h4557;
            4558: bcd <= 16'h4558;
            4559: bcd <= 16'h4559;
            4560: bcd <= 16'h4560;
            4561: bcd <= 16'h4561;
            4562: bcd <= 16'h4562;
            4563: bcd <= 16'h4563;
            4564: bcd <= 16'h4564;
            4565: bcd <= 16'h4565;
            4566: bcd <= 16'h4566;
            4567: bcd <= 16'h4567;
            4568: bcd <= 16'h4568;
            4569: bcd <= 16'h4569;
            4570: bcd <= 16'h4570;
            4571: bcd <= 16'h4571;
            4572: bcd <= 16'h4572;
            4573: bcd <= 16'h4573;
            4574: bcd <= 16'h4574;
            4575: bcd <= 16'h4575;
            4576: bcd <= 16'h4576;
            4577: bcd <= 16'h4577;
            4578: bcd <= 16'h4578;
            4579: bcd <= 16'h4579;
            4580: bcd <= 16'h4580;
            4581: bcd <= 16'h4581;
            4582: bcd <= 16'h4582;
            4583: bcd <= 16'h4583;
            4584: bcd <= 16'h4584;
            4585: bcd <= 16'h4585;
            4586: bcd <= 16'h4586;
            4587: bcd <= 16'h4587;
            4588: bcd <= 16'h4588;
            4589: bcd <= 16'h4589;
            4590: bcd <= 16'h4590;
            4591: bcd <= 16'h4591;
            4592: bcd <= 16'h4592;
            4593: bcd <= 16'h4593;
            4594: bcd <= 16'h4594;
            4595: bcd <= 16'h4595;
            4596: bcd <= 16'h4596;
            4597: bcd <= 16'h4597;
            4598: bcd <= 16'h4598;
            4599: bcd <= 16'h4599;
            4600: bcd <= 16'h4600;
            4601: bcd <= 16'h4601;
            4602: bcd <= 16'h4602;
            4603: bcd <= 16'h4603;
            4604: bcd <= 16'h4604;
            4605: bcd <= 16'h4605;
            4606: bcd <= 16'h4606;
            4607: bcd <= 16'h4607;
            4608: bcd <= 16'h4608;
            4609: bcd <= 16'h4609;
            4610: bcd <= 16'h4610;
            4611: bcd <= 16'h4611;
            4612: bcd <= 16'h4612;
            4613: bcd <= 16'h4613;
            4614: bcd <= 16'h4614;
            4615: bcd <= 16'h4615;
            4616: bcd <= 16'h4616;
            4617: bcd <= 16'h4617;
            4618: bcd <= 16'h4618;
            4619: bcd <= 16'h4619;
            4620: bcd <= 16'h4620;
            4621: bcd <= 16'h4621;
            4622: bcd <= 16'h4622;
            4623: bcd <= 16'h4623;
            4624: bcd <= 16'h4624;
            4625: bcd <= 16'h4625;
            4626: bcd <= 16'h4626;
            4627: bcd <= 16'h4627;
            4628: bcd <= 16'h4628;
            4629: bcd <= 16'h4629;
            4630: bcd <= 16'h4630;
            4631: bcd <= 16'h4631;
            4632: bcd <= 16'h4632;
            4633: bcd <= 16'h4633;
            4634: bcd <= 16'h4634;
            4635: bcd <= 16'h4635;
            4636: bcd <= 16'h4636;
            4637: bcd <= 16'h4637;
            4638: bcd <= 16'h4638;
            4639: bcd <= 16'h4639;
            4640: bcd <= 16'h4640;
            4641: bcd <= 16'h4641;
            4642: bcd <= 16'h4642;
            4643: bcd <= 16'h4643;
            4644: bcd <= 16'h4644;
            4645: bcd <= 16'h4645;
            4646: bcd <= 16'h4646;
            4647: bcd <= 16'h4647;
            4648: bcd <= 16'h4648;
            4649: bcd <= 16'h4649;
            4650: bcd <= 16'h4650;
            4651: bcd <= 16'h4651;
            4652: bcd <= 16'h4652;
            4653: bcd <= 16'h4653;
            4654: bcd <= 16'h4654;
            4655: bcd <= 16'h4655;
            4656: bcd <= 16'h4656;
            4657: bcd <= 16'h4657;
            4658: bcd <= 16'h4658;
            4659: bcd <= 16'h4659;
            4660: bcd <= 16'h4660;
            4661: bcd <= 16'h4661;
            4662: bcd <= 16'h4662;
            4663: bcd <= 16'h4663;
            4664: bcd <= 16'h4664;
            4665: bcd <= 16'h4665;
            4666: bcd <= 16'h4666;
            4667: bcd <= 16'h4667;
            4668: bcd <= 16'h4668;
            4669: bcd <= 16'h4669;
            4670: bcd <= 16'h4670;
            4671: bcd <= 16'h4671;
            4672: bcd <= 16'h4672;
            4673: bcd <= 16'h4673;
            4674: bcd <= 16'h4674;
            4675: bcd <= 16'h4675;
            4676: bcd <= 16'h4676;
            4677: bcd <= 16'h4677;
            4678: bcd <= 16'h4678;
            4679: bcd <= 16'h4679;
            4680: bcd <= 16'h4680;
            4681: bcd <= 16'h4681;
            4682: bcd <= 16'h4682;
            4683: bcd <= 16'h4683;
            4684: bcd <= 16'h4684;
            4685: bcd <= 16'h4685;
            4686: bcd <= 16'h4686;
            4687: bcd <= 16'h4687;
            4688: bcd <= 16'h4688;
            4689: bcd <= 16'h4689;
            4690: bcd <= 16'h4690;
            4691: bcd <= 16'h4691;
            4692: bcd <= 16'h4692;
            4693: bcd <= 16'h4693;
            4694: bcd <= 16'h4694;
            4695: bcd <= 16'h4695;
            4696: bcd <= 16'h4696;
            4697: bcd <= 16'h4697;
            4698: bcd <= 16'h4698;
            4699: bcd <= 16'h4699;
            4700: bcd <= 16'h4700;
            4701: bcd <= 16'h4701;
            4702: bcd <= 16'h4702;
            4703: bcd <= 16'h4703;
            4704: bcd <= 16'h4704;
            4705: bcd <= 16'h4705;
            4706: bcd <= 16'h4706;
            4707: bcd <= 16'h4707;
            4708: bcd <= 16'h4708;
            4709: bcd <= 16'h4709;
            4710: bcd <= 16'h4710;
            4711: bcd <= 16'h4711;
            4712: bcd <= 16'h4712;
            4713: bcd <= 16'h4713;
            4714: bcd <= 16'h4714;
            4715: bcd <= 16'h4715;
            4716: bcd <= 16'h4716;
            4717: bcd <= 16'h4717;
            4718: bcd <= 16'h4718;
            4719: bcd <= 16'h4719;
            4720: bcd <= 16'h4720;
            4721: bcd <= 16'h4721;
            4722: bcd <= 16'h4722;
            4723: bcd <= 16'h4723;
            4724: bcd <= 16'h4724;
            4725: bcd <= 16'h4725;
            4726: bcd <= 16'h4726;
            4727: bcd <= 16'h4727;
            4728: bcd <= 16'h4728;
            4729: bcd <= 16'h4729;
            4730: bcd <= 16'h4730;
            4731: bcd <= 16'h4731;
            4732: bcd <= 16'h4732;
            4733: bcd <= 16'h4733;
            4734: bcd <= 16'h4734;
            4735: bcd <= 16'h4735;
            4736: bcd <= 16'h4736;
            4737: bcd <= 16'h4737;
            4738: bcd <= 16'h4738;
            4739: bcd <= 16'h4739;
            4740: bcd <= 16'h4740;
            4741: bcd <= 16'h4741;
            4742: bcd <= 16'h4742;
            4743: bcd <= 16'h4743;
            4744: bcd <= 16'h4744;
            4745: bcd <= 16'h4745;
            4746: bcd <= 16'h4746;
            4747: bcd <= 16'h4747;
            4748: bcd <= 16'h4748;
            4749: bcd <= 16'h4749;
            4750: bcd <= 16'h4750;
            4751: bcd <= 16'h4751;
            4752: bcd <= 16'h4752;
            4753: bcd <= 16'h4753;
            4754: bcd <= 16'h4754;
            4755: bcd <= 16'h4755;
            4756: bcd <= 16'h4756;
            4757: bcd <= 16'h4757;
            4758: bcd <= 16'h4758;
            4759: bcd <= 16'h4759;
            4760: bcd <= 16'h4760;
            4761: bcd <= 16'h4761;
            4762: bcd <= 16'h4762;
            4763: bcd <= 16'h4763;
            4764: bcd <= 16'h4764;
            4765: bcd <= 16'h4765;
            4766: bcd <= 16'h4766;
            4767: bcd <= 16'h4767;
            4768: bcd <= 16'h4768;
            4769: bcd <= 16'h4769;
            4770: bcd <= 16'h4770;
            4771: bcd <= 16'h4771;
            4772: bcd <= 16'h4772;
            4773: bcd <= 16'h4773;
            4774: bcd <= 16'h4774;
            4775: bcd <= 16'h4775;
            4776: bcd <= 16'h4776;
            4777: bcd <= 16'h4777;
            4778: bcd <= 16'h4778;
            4779: bcd <= 16'h4779;
            4780: bcd <= 16'h4780;
            4781: bcd <= 16'h4781;
            4782: bcd <= 16'h4782;
            4783: bcd <= 16'h4783;
            4784: bcd <= 16'h4784;
            4785: bcd <= 16'h4785;
            4786: bcd <= 16'h4786;
            4787: bcd <= 16'h4787;
            4788: bcd <= 16'h4788;
            4789: bcd <= 16'h4789;
            4790: bcd <= 16'h4790;
            4791: bcd <= 16'h4791;
            4792: bcd <= 16'h4792;
            4793: bcd <= 16'h4793;
            4794: bcd <= 16'h4794;
            4795: bcd <= 16'h4795;
            4796: bcd <= 16'h4796;
            4797: bcd <= 16'h4797;
            4798: bcd <= 16'h4798;
            4799: bcd <= 16'h4799;
            4800: bcd <= 16'h4800;
            4801: bcd <= 16'h4801;
            4802: bcd <= 16'h4802;
            4803: bcd <= 16'h4803;
            4804: bcd <= 16'h4804;
            4805: bcd <= 16'h4805;
            4806: bcd <= 16'h4806;
            4807: bcd <= 16'h4807;
            4808: bcd <= 16'h4808;
            4809: bcd <= 16'h4809;
            4810: bcd <= 16'h4810;
            4811: bcd <= 16'h4811;
            4812: bcd <= 16'h4812;
            4813: bcd <= 16'h4813;
            4814: bcd <= 16'h4814;
            4815: bcd <= 16'h4815;
            4816: bcd <= 16'h4816;
            4817: bcd <= 16'h4817;
            4818: bcd <= 16'h4818;
            4819: bcd <= 16'h4819;
            4820: bcd <= 16'h4820;
            4821: bcd <= 16'h4821;
            4822: bcd <= 16'h4822;
            4823: bcd <= 16'h4823;
            4824: bcd <= 16'h4824;
            4825: bcd <= 16'h4825;
            4826: bcd <= 16'h4826;
            4827: bcd <= 16'h4827;
            4828: bcd <= 16'h4828;
            4829: bcd <= 16'h4829;
            4830: bcd <= 16'h4830;
            4831: bcd <= 16'h4831;
            4832: bcd <= 16'h4832;
            4833: bcd <= 16'h4833;
            4834: bcd <= 16'h4834;
            4835: bcd <= 16'h4835;
            4836: bcd <= 16'h4836;
            4837: bcd <= 16'h4837;
            4838: bcd <= 16'h4838;
            4839: bcd <= 16'h4839;
            4840: bcd <= 16'h4840;
            4841: bcd <= 16'h4841;
            4842: bcd <= 16'h4842;
            4843: bcd <= 16'h4843;
            4844: bcd <= 16'h4844;
            4845: bcd <= 16'h4845;
            4846: bcd <= 16'h4846;
            4847: bcd <= 16'h4847;
            4848: bcd <= 16'h4848;
            4849: bcd <= 16'h4849;
            4850: bcd <= 16'h4850;
            4851: bcd <= 16'h4851;
            4852: bcd <= 16'h4852;
            4853: bcd <= 16'h4853;
            4854: bcd <= 16'h4854;
            4855: bcd <= 16'h4855;
            4856: bcd <= 16'h4856;
            4857: bcd <= 16'h4857;
            4858: bcd <= 16'h4858;
            4859: bcd <= 16'h4859;
            4860: bcd <= 16'h4860;
            4861: bcd <= 16'h4861;
            4862: bcd <= 16'h4862;
            4863: bcd <= 16'h4863;
            4864: bcd <= 16'h4864;
            4865: bcd <= 16'h4865;
            4866: bcd <= 16'h4866;
            4867: bcd <= 16'h4867;
            4868: bcd <= 16'h4868;
            4869: bcd <= 16'h4869;
            4870: bcd <= 16'h4870;
            4871: bcd <= 16'h4871;
            4872: bcd <= 16'h4872;
            4873: bcd <= 16'h4873;
            4874: bcd <= 16'h4874;
            4875: bcd <= 16'h4875;
            4876: bcd <= 16'h4876;
            4877: bcd <= 16'h4877;
            4878: bcd <= 16'h4878;
            4879: bcd <= 16'h4879;
            4880: bcd <= 16'h4880;
            4881: bcd <= 16'h4881;
            4882: bcd <= 16'h4882;
            4883: bcd <= 16'h4883;
            4884: bcd <= 16'h4884;
            4885: bcd <= 16'h4885;
            4886: bcd <= 16'h4886;
            4887: bcd <= 16'h4887;
            4888: bcd <= 16'h4888;
            4889: bcd <= 16'h4889;
            4890: bcd <= 16'h4890;
            4891: bcd <= 16'h4891;
            4892: bcd <= 16'h4892;
            4893: bcd <= 16'h4893;
            4894: bcd <= 16'h4894;
            4895: bcd <= 16'h4895;
            4896: bcd <= 16'h4896;
            4897: bcd <= 16'h4897;
            4898: bcd <= 16'h4898;
            4899: bcd <= 16'h4899;
            4900: bcd <= 16'h4900;
            4901: bcd <= 16'h4901;
            4902: bcd <= 16'h4902;
            4903: bcd <= 16'h4903;
            4904: bcd <= 16'h4904;
            4905: bcd <= 16'h4905;
            4906: bcd <= 16'h4906;
            4907: bcd <= 16'h4907;
            4908: bcd <= 16'h4908;
            4909: bcd <= 16'h4909;
            4910: bcd <= 16'h4910;
            4911: bcd <= 16'h4911;
            4912: bcd <= 16'h4912;
            4913: bcd <= 16'h4913;
            4914: bcd <= 16'h4914;
            4915: bcd <= 16'h4915;
            4916: bcd <= 16'h4916;
            4917: bcd <= 16'h4917;
            4918: bcd <= 16'h4918;
            4919: bcd <= 16'h4919;
            4920: bcd <= 16'h4920;
            4921: bcd <= 16'h4921;
            4922: bcd <= 16'h4922;
            4923: bcd <= 16'h4923;
            4924: bcd <= 16'h4924;
            4925: bcd <= 16'h4925;
            4926: bcd <= 16'h4926;
            4927: bcd <= 16'h4927;
            4928: bcd <= 16'h4928;
            4929: bcd <= 16'h4929;
            4930: bcd <= 16'h4930;
            4931: bcd <= 16'h4931;
            4932: bcd <= 16'h4932;
            4933: bcd <= 16'h4933;
            4934: bcd <= 16'h4934;
            4935: bcd <= 16'h4935;
            4936: bcd <= 16'h4936;
            4937: bcd <= 16'h4937;
            4938: bcd <= 16'h4938;
            4939: bcd <= 16'h4939;
            4940: bcd <= 16'h4940;
            4941: bcd <= 16'h4941;
            4942: bcd <= 16'h4942;
            4943: bcd <= 16'h4943;
            4944: bcd <= 16'h4944;
            4945: bcd <= 16'h4945;
            4946: bcd <= 16'h4946;
            4947: bcd <= 16'h4947;
            4948: bcd <= 16'h4948;
            4949: bcd <= 16'h4949;
            4950: bcd <= 16'h4950;
            4951: bcd <= 16'h4951;
            4952: bcd <= 16'h4952;
            4953: bcd <= 16'h4953;
            4954: bcd <= 16'h4954;
            4955: bcd <= 16'h4955;
            4956: bcd <= 16'h4956;
            4957: bcd <= 16'h4957;
            4958: bcd <= 16'h4958;
            4959: bcd <= 16'h4959;
            4960: bcd <= 16'h4960;
            4961: bcd <= 16'h4961;
            4962: bcd <= 16'h4962;
            4963: bcd <= 16'h4963;
            4964: bcd <= 16'h4964;
            4965: bcd <= 16'h4965;
            4966: bcd <= 16'h4966;
            4967: bcd <= 16'h4967;
            4968: bcd <= 16'h4968;
            4969: bcd <= 16'h4969;
            4970: bcd <= 16'h4970;
            4971: bcd <= 16'h4971;
            4972: bcd <= 16'h4972;
            4973: bcd <= 16'h4973;
            4974: bcd <= 16'h4974;
            4975: bcd <= 16'h4975;
            4976: bcd <= 16'h4976;
            4977: bcd <= 16'h4977;
            4978: bcd <= 16'h4978;
            4979: bcd <= 16'h4979;
            4980: bcd <= 16'h4980;
            4981: bcd <= 16'h4981;
            4982: bcd <= 16'h4982;
            4983: bcd <= 16'h4983;
            4984: bcd <= 16'h4984;
            4985: bcd <= 16'h4985;
            4986: bcd <= 16'h4986;
            4987: bcd <= 16'h4987;
            4988: bcd <= 16'h4988;
            4989: bcd <= 16'h4989;
            4990: bcd <= 16'h4990;
            4991: bcd <= 16'h4991;
            4992: bcd <= 16'h4992;
            4993: bcd <= 16'h4993;
            4994: bcd <= 16'h4994;
            4995: bcd <= 16'h4995;
            4996: bcd <= 16'h4996;
            4997: bcd <= 16'h4997;
            4998: bcd <= 16'h4998;
            4999: bcd <= 16'h4999;
            5000: bcd <= 16'h5000;
            5001: bcd <= 16'h5001;
            5002: bcd <= 16'h5002;
            5003: bcd <= 16'h5003;
            5004: bcd <= 16'h5004;
            5005: bcd <= 16'h5005;
            5006: bcd <= 16'h5006;
            5007: bcd <= 16'h5007;
            5008: bcd <= 16'h5008;
            5009: bcd <= 16'h5009;
            5010: bcd <= 16'h5010;
            5011: bcd <= 16'h5011;
            5012: bcd <= 16'h5012;
            5013: bcd <= 16'h5013;
            5014: bcd <= 16'h5014;
            5015: bcd <= 16'h5015;
            5016: bcd <= 16'h5016;
            5017: bcd <= 16'h5017;
            5018: bcd <= 16'h5018;
            5019: bcd <= 16'h5019;
            5020: bcd <= 16'h5020;
            5021: bcd <= 16'h5021;
            5022: bcd <= 16'h5022;
            5023: bcd <= 16'h5023;
            5024: bcd <= 16'h5024;
            5025: bcd <= 16'h5025;
            5026: bcd <= 16'h5026;
            5027: bcd <= 16'h5027;
            5028: bcd <= 16'h5028;
            5029: bcd <= 16'h5029;
            5030: bcd <= 16'h5030;
            5031: bcd <= 16'h5031;
            5032: bcd <= 16'h5032;
            5033: bcd <= 16'h5033;
            5034: bcd <= 16'h5034;
            5035: bcd <= 16'h5035;
            5036: bcd <= 16'h5036;
            5037: bcd <= 16'h5037;
            5038: bcd <= 16'h5038;
            5039: bcd <= 16'h5039;
            5040: bcd <= 16'h5040;
            5041: bcd <= 16'h5041;
            5042: bcd <= 16'h5042;
            5043: bcd <= 16'h5043;
            5044: bcd <= 16'h5044;
            5045: bcd <= 16'h5045;
            5046: bcd <= 16'h5046;
            5047: bcd <= 16'h5047;
            5048: bcd <= 16'h5048;
            5049: bcd <= 16'h5049;
            5050: bcd <= 16'h5050;
            5051: bcd <= 16'h5051;
            5052: bcd <= 16'h5052;
            5053: bcd <= 16'h5053;
            5054: bcd <= 16'h5054;
            5055: bcd <= 16'h5055;
            5056: bcd <= 16'h5056;
            5057: bcd <= 16'h5057;
            5058: bcd <= 16'h5058;
            5059: bcd <= 16'h5059;
            5060: bcd <= 16'h5060;
            5061: bcd <= 16'h5061;
            5062: bcd <= 16'h5062;
            5063: bcd <= 16'h5063;
            5064: bcd <= 16'h5064;
            5065: bcd <= 16'h5065;
            5066: bcd <= 16'h5066;
            5067: bcd <= 16'h5067;
            5068: bcd <= 16'h5068;
            5069: bcd <= 16'h5069;
            5070: bcd <= 16'h5070;
            5071: bcd <= 16'h5071;
            5072: bcd <= 16'h5072;
            5073: bcd <= 16'h5073;
            5074: bcd <= 16'h5074;
            5075: bcd <= 16'h5075;
            5076: bcd <= 16'h5076;
            5077: bcd <= 16'h5077;
            5078: bcd <= 16'h5078;
            5079: bcd <= 16'h5079;
            5080: bcd <= 16'h5080;
            5081: bcd <= 16'h5081;
            5082: bcd <= 16'h5082;
            5083: bcd <= 16'h5083;
            5084: bcd <= 16'h5084;
            5085: bcd <= 16'h5085;
            5086: bcd <= 16'h5086;
            5087: bcd <= 16'h5087;
            5088: bcd <= 16'h5088;
            5089: bcd <= 16'h5089;
            5090: bcd <= 16'h5090;
            5091: bcd <= 16'h5091;
            5092: bcd <= 16'h5092;
            5093: bcd <= 16'h5093;
            5094: bcd <= 16'h5094;
            5095: bcd <= 16'h5095;
            5096: bcd <= 16'h5096;
            5097: bcd <= 16'h5097;
            5098: bcd <= 16'h5098;
            5099: bcd <= 16'h5099;
            5100: bcd <= 16'h5100;
            5101: bcd <= 16'h5101;
            5102: bcd <= 16'h5102;
            5103: bcd <= 16'h5103;
            5104: bcd <= 16'h5104;
            5105: bcd <= 16'h5105;
            5106: bcd <= 16'h5106;
            5107: bcd <= 16'h5107;
            5108: bcd <= 16'h5108;
            5109: bcd <= 16'h5109;
            5110: bcd <= 16'h5110;
            5111: bcd <= 16'h5111;
            5112: bcd <= 16'h5112;
            5113: bcd <= 16'h5113;
            5114: bcd <= 16'h5114;
            5115: bcd <= 16'h5115;
            5116: bcd <= 16'h5116;
            5117: bcd <= 16'h5117;
            5118: bcd <= 16'h5118;
            5119: bcd <= 16'h5119;
            5120: bcd <= 16'h5120;
            5121: bcd <= 16'h5121;
            5122: bcd <= 16'h5122;
            5123: bcd <= 16'h5123;
            5124: bcd <= 16'h5124;
            5125: bcd <= 16'h5125;
            5126: bcd <= 16'h5126;
            5127: bcd <= 16'h5127;
            5128: bcd <= 16'h5128;
            5129: bcd <= 16'h5129;
            5130: bcd <= 16'h5130;
            5131: bcd <= 16'h5131;
            5132: bcd <= 16'h5132;
            5133: bcd <= 16'h5133;
            5134: bcd <= 16'h5134;
            5135: bcd <= 16'h5135;
            5136: bcd <= 16'h5136;
            5137: bcd <= 16'h5137;
            5138: bcd <= 16'h5138;
            5139: bcd <= 16'h5139;
            5140: bcd <= 16'h5140;
            5141: bcd <= 16'h5141;
            5142: bcd <= 16'h5142;
            5143: bcd <= 16'h5143;
            5144: bcd <= 16'h5144;
            5145: bcd <= 16'h5145;
            5146: bcd <= 16'h5146;
            5147: bcd <= 16'h5147;
            5148: bcd <= 16'h5148;
            5149: bcd <= 16'h5149;
            5150: bcd <= 16'h5150;
            5151: bcd <= 16'h5151;
            5152: bcd <= 16'h5152;
            5153: bcd <= 16'h5153;
            5154: bcd <= 16'h5154;
            5155: bcd <= 16'h5155;
            5156: bcd <= 16'h5156;
            5157: bcd <= 16'h5157;
            5158: bcd <= 16'h5158;
            5159: bcd <= 16'h5159;
            5160: bcd <= 16'h5160;
            5161: bcd <= 16'h5161;
            5162: bcd <= 16'h5162;
            5163: bcd <= 16'h5163;
            5164: bcd <= 16'h5164;
            5165: bcd <= 16'h5165;
            5166: bcd <= 16'h5166;
            5167: bcd <= 16'h5167;
            5168: bcd <= 16'h5168;
            5169: bcd <= 16'h5169;
            5170: bcd <= 16'h5170;
            5171: bcd <= 16'h5171;
            5172: bcd <= 16'h5172;
            5173: bcd <= 16'h5173;
            5174: bcd <= 16'h5174;
            5175: bcd <= 16'h5175;
            5176: bcd <= 16'h5176;
            5177: bcd <= 16'h5177;
            5178: bcd <= 16'h5178;
            5179: bcd <= 16'h5179;
            5180: bcd <= 16'h5180;
            5181: bcd <= 16'h5181;
            5182: bcd <= 16'h5182;
            5183: bcd <= 16'h5183;
            5184: bcd <= 16'h5184;
            5185: bcd <= 16'h5185;
            5186: bcd <= 16'h5186;
            5187: bcd <= 16'h5187;
            5188: bcd <= 16'h5188;
            5189: bcd <= 16'h5189;
            5190: bcd <= 16'h5190;
            5191: bcd <= 16'h5191;
            5192: bcd <= 16'h5192;
            5193: bcd <= 16'h5193;
            5194: bcd <= 16'h5194;
            5195: bcd <= 16'h5195;
            5196: bcd <= 16'h5196;
            5197: bcd <= 16'h5197;
            5198: bcd <= 16'h5198;
            5199: bcd <= 16'h5199;
            5200: bcd <= 16'h5200;
            5201: bcd <= 16'h5201;
            5202: bcd <= 16'h5202;
            5203: bcd <= 16'h5203;
            5204: bcd <= 16'h5204;
            5205: bcd <= 16'h5205;
            5206: bcd <= 16'h5206;
            5207: bcd <= 16'h5207;
            5208: bcd <= 16'h5208;
            5209: bcd <= 16'h5209;
            5210: bcd <= 16'h5210;
            5211: bcd <= 16'h5211;
            5212: bcd <= 16'h5212;
            5213: bcd <= 16'h5213;
            5214: bcd <= 16'h5214;
            5215: bcd <= 16'h5215;
            5216: bcd <= 16'h5216;
            5217: bcd <= 16'h5217;
            5218: bcd <= 16'h5218;
            5219: bcd <= 16'h5219;
            5220: bcd <= 16'h5220;
            5221: bcd <= 16'h5221;
            5222: bcd <= 16'h5222;
            5223: bcd <= 16'h5223;
            5224: bcd <= 16'h5224;
            5225: bcd <= 16'h5225;
            5226: bcd <= 16'h5226;
            5227: bcd <= 16'h5227;
            5228: bcd <= 16'h5228;
            5229: bcd <= 16'h5229;
            5230: bcd <= 16'h5230;
            5231: bcd <= 16'h5231;
            5232: bcd <= 16'h5232;
            5233: bcd <= 16'h5233;
            5234: bcd <= 16'h5234;
            5235: bcd <= 16'h5235;
            5236: bcd <= 16'h5236;
            5237: bcd <= 16'h5237;
            5238: bcd <= 16'h5238;
            5239: bcd <= 16'h5239;
            5240: bcd <= 16'h5240;
            5241: bcd <= 16'h5241;
            5242: bcd <= 16'h5242;
            5243: bcd <= 16'h5243;
            5244: bcd <= 16'h5244;
            5245: bcd <= 16'h5245;
            5246: bcd <= 16'h5246;
            5247: bcd <= 16'h5247;
            5248: bcd <= 16'h5248;
            5249: bcd <= 16'h5249;
            5250: bcd <= 16'h5250;
            5251: bcd <= 16'h5251;
            5252: bcd <= 16'h5252;
            5253: bcd <= 16'h5253;
            5254: bcd <= 16'h5254;
            5255: bcd <= 16'h5255;
            5256: bcd <= 16'h5256;
            5257: bcd <= 16'h5257;
            5258: bcd <= 16'h5258;
            5259: bcd <= 16'h5259;
            5260: bcd <= 16'h5260;
            5261: bcd <= 16'h5261;
            5262: bcd <= 16'h5262;
            5263: bcd <= 16'h5263;
            5264: bcd <= 16'h5264;
            5265: bcd <= 16'h5265;
            5266: bcd <= 16'h5266;
            5267: bcd <= 16'h5267;
            5268: bcd <= 16'h5268;
            5269: bcd <= 16'h5269;
            5270: bcd <= 16'h5270;
            5271: bcd <= 16'h5271;
            5272: bcd <= 16'h5272;
            5273: bcd <= 16'h5273;
            5274: bcd <= 16'h5274;
            5275: bcd <= 16'h5275;
            5276: bcd <= 16'h5276;
            5277: bcd <= 16'h5277;
            5278: bcd <= 16'h5278;
            5279: bcd <= 16'h5279;
            5280: bcd <= 16'h5280;
            5281: bcd <= 16'h5281;
            5282: bcd <= 16'h5282;
            5283: bcd <= 16'h5283;
            5284: bcd <= 16'h5284;
            5285: bcd <= 16'h5285;
            5286: bcd <= 16'h5286;
            5287: bcd <= 16'h5287;
            5288: bcd <= 16'h5288;
            5289: bcd <= 16'h5289;
            5290: bcd <= 16'h5290;
            5291: bcd <= 16'h5291;
            5292: bcd <= 16'h5292;
            5293: bcd <= 16'h5293;
            5294: bcd <= 16'h5294;
            5295: bcd <= 16'h5295;
            5296: bcd <= 16'h5296;
            5297: bcd <= 16'h5297;
            5298: bcd <= 16'h5298;
            5299: bcd <= 16'h5299;
            5300: bcd <= 16'h5300;
            5301: bcd <= 16'h5301;
            5302: bcd <= 16'h5302;
            5303: bcd <= 16'h5303;
            5304: bcd <= 16'h5304;
            5305: bcd <= 16'h5305;
            5306: bcd <= 16'h5306;
            5307: bcd <= 16'h5307;
            5308: bcd <= 16'h5308;
            5309: bcd <= 16'h5309;
            5310: bcd <= 16'h5310;
            5311: bcd <= 16'h5311;
            5312: bcd <= 16'h5312;
            5313: bcd <= 16'h5313;
            5314: bcd <= 16'h5314;
            5315: bcd <= 16'h5315;
            5316: bcd <= 16'h5316;
            5317: bcd <= 16'h5317;
            5318: bcd <= 16'h5318;
            5319: bcd <= 16'h5319;
            5320: bcd <= 16'h5320;
            5321: bcd <= 16'h5321;
            5322: bcd <= 16'h5322;
            5323: bcd <= 16'h5323;
            5324: bcd <= 16'h5324;
            5325: bcd <= 16'h5325;
            5326: bcd <= 16'h5326;
            5327: bcd <= 16'h5327;
            5328: bcd <= 16'h5328;
            5329: bcd <= 16'h5329;
            5330: bcd <= 16'h5330;
            5331: bcd <= 16'h5331;
            5332: bcd <= 16'h5332;
            5333: bcd <= 16'h5333;
            5334: bcd <= 16'h5334;
            5335: bcd <= 16'h5335;
            5336: bcd <= 16'h5336;
            5337: bcd <= 16'h5337;
            5338: bcd <= 16'h5338;
            5339: bcd <= 16'h5339;
            5340: bcd <= 16'h5340;
            5341: bcd <= 16'h5341;
            5342: bcd <= 16'h5342;
            5343: bcd <= 16'h5343;
            5344: bcd <= 16'h5344;
            5345: bcd <= 16'h5345;
            5346: bcd <= 16'h5346;
            5347: bcd <= 16'h5347;
            5348: bcd <= 16'h5348;
            5349: bcd <= 16'h5349;
            5350: bcd <= 16'h5350;
            5351: bcd <= 16'h5351;
            5352: bcd <= 16'h5352;
            5353: bcd <= 16'h5353;
            5354: bcd <= 16'h5354;
            5355: bcd <= 16'h5355;
            5356: bcd <= 16'h5356;
            5357: bcd <= 16'h5357;
            5358: bcd <= 16'h5358;
            5359: bcd <= 16'h5359;
            5360: bcd <= 16'h5360;
            5361: bcd <= 16'h5361;
            5362: bcd <= 16'h5362;
            5363: bcd <= 16'h5363;
            5364: bcd <= 16'h5364;
            5365: bcd <= 16'h5365;
            5366: bcd <= 16'h5366;
            5367: bcd <= 16'h5367;
            5368: bcd <= 16'h5368;
            5369: bcd <= 16'h5369;
            5370: bcd <= 16'h5370;
            5371: bcd <= 16'h5371;
            5372: bcd <= 16'h5372;
            5373: bcd <= 16'h5373;
            5374: bcd <= 16'h5374;
            5375: bcd <= 16'h5375;
            5376: bcd <= 16'h5376;
            5377: bcd <= 16'h5377;
            5378: bcd <= 16'h5378;
            5379: bcd <= 16'h5379;
            5380: bcd <= 16'h5380;
            5381: bcd <= 16'h5381;
            5382: bcd <= 16'h5382;
            5383: bcd <= 16'h5383;
            5384: bcd <= 16'h5384;
            5385: bcd <= 16'h5385;
            5386: bcd <= 16'h5386;
            5387: bcd <= 16'h5387;
            5388: bcd <= 16'h5388;
            5389: bcd <= 16'h5389;
            5390: bcd <= 16'h5390;
            5391: bcd <= 16'h5391;
            5392: bcd <= 16'h5392;
            5393: bcd <= 16'h5393;
            5394: bcd <= 16'h5394;
            5395: bcd <= 16'h5395;
            5396: bcd <= 16'h5396;
            5397: bcd <= 16'h5397;
            5398: bcd <= 16'h5398;
            5399: bcd <= 16'h5399;
            5400: bcd <= 16'h5400;
            5401: bcd <= 16'h5401;
            5402: bcd <= 16'h5402;
            5403: bcd <= 16'h5403;
            5404: bcd <= 16'h5404;
            5405: bcd <= 16'h5405;
            5406: bcd <= 16'h5406;
            5407: bcd <= 16'h5407;
            5408: bcd <= 16'h5408;
            5409: bcd <= 16'h5409;
            5410: bcd <= 16'h5410;
            5411: bcd <= 16'h5411;
            5412: bcd <= 16'h5412;
            5413: bcd <= 16'h5413;
            5414: bcd <= 16'h5414;
            5415: bcd <= 16'h5415;
            5416: bcd <= 16'h5416;
            5417: bcd <= 16'h5417;
            5418: bcd <= 16'h5418;
            5419: bcd <= 16'h5419;
            5420: bcd <= 16'h5420;
            5421: bcd <= 16'h5421;
            5422: bcd <= 16'h5422;
            5423: bcd <= 16'h5423;
            5424: bcd <= 16'h5424;
            5425: bcd <= 16'h5425;
            5426: bcd <= 16'h5426;
            5427: bcd <= 16'h5427;
            5428: bcd <= 16'h5428;
            5429: bcd <= 16'h5429;
            5430: bcd <= 16'h5430;
            5431: bcd <= 16'h5431;
            5432: bcd <= 16'h5432;
            5433: bcd <= 16'h5433;
            5434: bcd <= 16'h5434;
            5435: bcd <= 16'h5435;
            5436: bcd <= 16'h5436;
            5437: bcd <= 16'h5437;
            5438: bcd <= 16'h5438;
            5439: bcd <= 16'h5439;
            5440: bcd <= 16'h5440;
            5441: bcd <= 16'h5441;
            5442: bcd <= 16'h5442;
            5443: bcd <= 16'h5443;
            5444: bcd <= 16'h5444;
            5445: bcd <= 16'h5445;
            5446: bcd <= 16'h5446;
            5447: bcd <= 16'h5447;
            5448: bcd <= 16'h5448;
            5449: bcd <= 16'h5449;
            5450: bcd <= 16'h5450;
            5451: bcd <= 16'h5451;
            5452: bcd <= 16'h5452;
            5453: bcd <= 16'h5453;
            5454: bcd <= 16'h5454;
            5455: bcd <= 16'h5455;
            5456: bcd <= 16'h5456;
            5457: bcd <= 16'h5457;
            5458: bcd <= 16'h5458;
            5459: bcd <= 16'h5459;
            5460: bcd <= 16'h5460;
            5461: bcd <= 16'h5461;
            5462: bcd <= 16'h5462;
            5463: bcd <= 16'h5463;
            5464: bcd <= 16'h5464;
            5465: bcd <= 16'h5465;
            5466: bcd <= 16'h5466;
            5467: bcd <= 16'h5467;
            5468: bcd <= 16'h5468;
            5469: bcd <= 16'h5469;
            5470: bcd <= 16'h5470;
            5471: bcd <= 16'h5471;
            5472: bcd <= 16'h5472;
            5473: bcd <= 16'h5473;
            5474: bcd <= 16'h5474;
            5475: bcd <= 16'h5475;
            5476: bcd <= 16'h5476;
            5477: bcd <= 16'h5477;
            5478: bcd <= 16'h5478;
            5479: bcd <= 16'h5479;
            5480: bcd <= 16'h5480;
            5481: bcd <= 16'h5481;
            5482: bcd <= 16'h5482;
            5483: bcd <= 16'h5483;
            5484: bcd <= 16'h5484;
            5485: bcd <= 16'h5485;
            5486: bcd <= 16'h5486;
            5487: bcd <= 16'h5487;
            5488: bcd <= 16'h5488;
            5489: bcd <= 16'h5489;
            5490: bcd <= 16'h5490;
            5491: bcd <= 16'h5491;
            5492: bcd <= 16'h5492;
            5493: bcd <= 16'h5493;
            5494: bcd <= 16'h5494;
            5495: bcd <= 16'h5495;
            5496: bcd <= 16'h5496;
            5497: bcd <= 16'h5497;
            5498: bcd <= 16'h5498;
            5499: bcd <= 16'h5499;
            5500: bcd <= 16'h5500;
            5501: bcd <= 16'h5501;
            5502: bcd <= 16'h5502;
            5503: bcd <= 16'h5503;
            5504: bcd <= 16'h5504;
            5505: bcd <= 16'h5505;
            5506: bcd <= 16'h5506;
            5507: bcd <= 16'h5507;
            5508: bcd <= 16'h5508;
            5509: bcd <= 16'h5509;
            5510: bcd <= 16'h5510;
            5511: bcd <= 16'h5511;
            5512: bcd <= 16'h5512;
            5513: bcd <= 16'h5513;
            5514: bcd <= 16'h5514;
            5515: bcd <= 16'h5515;
            5516: bcd <= 16'h5516;
            5517: bcd <= 16'h5517;
            5518: bcd <= 16'h5518;
            5519: bcd <= 16'h5519;
            5520: bcd <= 16'h5520;
            5521: bcd <= 16'h5521;
            5522: bcd <= 16'h5522;
            5523: bcd <= 16'h5523;
            5524: bcd <= 16'h5524;
            5525: bcd <= 16'h5525;
            5526: bcd <= 16'h5526;
            5527: bcd <= 16'h5527;
            5528: bcd <= 16'h5528;
            5529: bcd <= 16'h5529;
            5530: bcd <= 16'h5530;
            5531: bcd <= 16'h5531;
            5532: bcd <= 16'h5532;
            5533: bcd <= 16'h5533;
            5534: bcd <= 16'h5534;
            5535: bcd <= 16'h5535;
            5536: bcd <= 16'h5536;
            5537: bcd <= 16'h5537;
            5538: bcd <= 16'h5538;
            5539: bcd <= 16'h5539;
            5540: bcd <= 16'h5540;
            5541: bcd <= 16'h5541;
            5542: bcd <= 16'h5542;
            5543: bcd <= 16'h5543;
            5544: bcd <= 16'h5544;
            5545: bcd <= 16'h5545;
            5546: bcd <= 16'h5546;
            5547: bcd <= 16'h5547;
            5548: bcd <= 16'h5548;
            5549: bcd <= 16'h5549;
            5550: bcd <= 16'h5550;
            5551: bcd <= 16'h5551;
            5552: bcd <= 16'h5552;
            5553: bcd <= 16'h5553;
            5554: bcd <= 16'h5554;
            5555: bcd <= 16'h5555;
            5556: bcd <= 16'h5556;
            5557: bcd <= 16'h5557;
            5558: bcd <= 16'h5558;
            5559: bcd <= 16'h5559;
            5560: bcd <= 16'h5560;
            5561: bcd <= 16'h5561;
            5562: bcd <= 16'h5562;
            5563: bcd <= 16'h5563;
            5564: bcd <= 16'h5564;
            5565: bcd <= 16'h5565;
            5566: bcd <= 16'h5566;
            5567: bcd <= 16'h5567;
            5568: bcd <= 16'h5568;
            5569: bcd <= 16'h5569;
            5570: bcd <= 16'h5570;
            5571: bcd <= 16'h5571;
            5572: bcd <= 16'h5572;
            5573: bcd <= 16'h5573;
            5574: bcd <= 16'h5574;
            5575: bcd <= 16'h5575;
            5576: bcd <= 16'h5576;
            5577: bcd <= 16'h5577;
            5578: bcd <= 16'h5578;
            5579: bcd <= 16'h5579;
            5580: bcd <= 16'h5580;
            5581: bcd <= 16'h5581;
            5582: bcd <= 16'h5582;
            5583: bcd <= 16'h5583;
            5584: bcd <= 16'h5584;
            5585: bcd <= 16'h5585;
            5586: bcd <= 16'h5586;
            5587: bcd <= 16'h5587;
            5588: bcd <= 16'h5588;
            5589: bcd <= 16'h5589;
            5590: bcd <= 16'h5590;
            5591: bcd <= 16'h5591;
            5592: bcd <= 16'h5592;
            5593: bcd <= 16'h5593;
            5594: bcd <= 16'h5594;
            5595: bcd <= 16'h5595;
            5596: bcd <= 16'h5596;
            5597: bcd <= 16'h5597;
            5598: bcd <= 16'h5598;
            5599: bcd <= 16'h5599;
            5600: bcd <= 16'h5600;
            5601: bcd <= 16'h5601;
            5602: bcd <= 16'h5602;
            5603: bcd <= 16'h5603;
            5604: bcd <= 16'h5604;
            5605: bcd <= 16'h5605;
            5606: bcd <= 16'h5606;
            5607: bcd <= 16'h5607;
            5608: bcd <= 16'h5608;
            5609: bcd <= 16'h5609;
            5610: bcd <= 16'h5610;
            5611: bcd <= 16'h5611;
            5612: bcd <= 16'h5612;
            5613: bcd <= 16'h5613;
            5614: bcd <= 16'h5614;
            5615: bcd <= 16'h5615;
            5616: bcd <= 16'h5616;
            5617: bcd <= 16'h5617;
            5618: bcd <= 16'h5618;
            5619: bcd <= 16'h5619;
            5620: bcd <= 16'h5620;
            5621: bcd <= 16'h5621;
            5622: bcd <= 16'h5622;
            5623: bcd <= 16'h5623;
            5624: bcd <= 16'h5624;
            5625: bcd <= 16'h5625;
            5626: bcd <= 16'h5626;
            5627: bcd <= 16'h5627;
            5628: bcd <= 16'h5628;
            5629: bcd <= 16'h5629;
            5630: bcd <= 16'h5630;
            5631: bcd <= 16'h5631;
            5632: bcd <= 16'h5632;
            5633: bcd <= 16'h5633;
            5634: bcd <= 16'h5634;
            5635: bcd <= 16'h5635;
            5636: bcd <= 16'h5636;
            5637: bcd <= 16'h5637;
            5638: bcd <= 16'h5638;
            5639: bcd <= 16'h5639;
            5640: bcd <= 16'h5640;
            5641: bcd <= 16'h5641;
            5642: bcd <= 16'h5642;
            5643: bcd <= 16'h5643;
            5644: bcd <= 16'h5644;
            5645: bcd <= 16'h5645;
            5646: bcd <= 16'h5646;
            5647: bcd <= 16'h5647;
            5648: bcd <= 16'h5648;
            5649: bcd <= 16'h5649;
            5650: bcd <= 16'h5650;
            5651: bcd <= 16'h5651;
            5652: bcd <= 16'h5652;
            5653: bcd <= 16'h5653;
            5654: bcd <= 16'h5654;
            5655: bcd <= 16'h5655;
            5656: bcd <= 16'h5656;
            5657: bcd <= 16'h5657;
            5658: bcd <= 16'h5658;
            5659: bcd <= 16'h5659;
            5660: bcd <= 16'h5660;
            5661: bcd <= 16'h5661;
            5662: bcd <= 16'h5662;
            5663: bcd <= 16'h5663;
            5664: bcd <= 16'h5664;
            5665: bcd <= 16'h5665;
            5666: bcd <= 16'h5666;
            5667: bcd <= 16'h5667;
            5668: bcd <= 16'h5668;
            5669: bcd <= 16'h5669;
            5670: bcd <= 16'h5670;
            5671: bcd <= 16'h5671;
            5672: bcd <= 16'h5672;
            5673: bcd <= 16'h5673;
            5674: bcd <= 16'h5674;
            5675: bcd <= 16'h5675;
            5676: bcd <= 16'h5676;
            5677: bcd <= 16'h5677;
            5678: bcd <= 16'h5678;
            5679: bcd <= 16'h5679;
            5680: bcd <= 16'h5680;
            5681: bcd <= 16'h5681;
            5682: bcd <= 16'h5682;
            5683: bcd <= 16'h5683;
            5684: bcd <= 16'h5684;
            5685: bcd <= 16'h5685;
            5686: bcd <= 16'h5686;
            5687: bcd <= 16'h5687;
            5688: bcd <= 16'h5688;
            5689: bcd <= 16'h5689;
            5690: bcd <= 16'h5690;
            5691: bcd <= 16'h5691;
            5692: bcd <= 16'h5692;
            5693: bcd <= 16'h5693;
            5694: bcd <= 16'h5694;
            5695: bcd <= 16'h5695;
            5696: bcd <= 16'h5696;
            5697: bcd <= 16'h5697;
            5698: bcd <= 16'h5698;
            5699: bcd <= 16'h5699;
            5700: bcd <= 16'h5700;
            5701: bcd <= 16'h5701;
            5702: bcd <= 16'h5702;
            5703: bcd <= 16'h5703;
            5704: bcd <= 16'h5704;
            5705: bcd <= 16'h5705;
            5706: bcd <= 16'h5706;
            5707: bcd <= 16'h5707;
            5708: bcd <= 16'h5708;
            5709: bcd <= 16'h5709;
            5710: bcd <= 16'h5710;
            5711: bcd <= 16'h5711;
            5712: bcd <= 16'h5712;
            5713: bcd <= 16'h5713;
            5714: bcd <= 16'h5714;
            5715: bcd <= 16'h5715;
            5716: bcd <= 16'h5716;
            5717: bcd <= 16'h5717;
            5718: bcd <= 16'h5718;
            5719: bcd <= 16'h5719;
            5720: bcd <= 16'h5720;
            5721: bcd <= 16'h5721;
            5722: bcd <= 16'h5722;
            5723: bcd <= 16'h5723;
            5724: bcd <= 16'h5724;
            5725: bcd <= 16'h5725;
            5726: bcd <= 16'h5726;
            5727: bcd <= 16'h5727;
            5728: bcd <= 16'h5728;
            5729: bcd <= 16'h5729;
            5730: bcd <= 16'h5730;
            5731: bcd <= 16'h5731;
            5732: bcd <= 16'h5732;
            5733: bcd <= 16'h5733;
            5734: bcd <= 16'h5734;
            5735: bcd <= 16'h5735;
            5736: bcd <= 16'h5736;
            5737: bcd <= 16'h5737;
            5738: bcd <= 16'h5738;
            5739: bcd <= 16'h5739;
            5740: bcd <= 16'h5740;
            5741: bcd <= 16'h5741;
            5742: bcd <= 16'h5742;
            5743: bcd <= 16'h5743;
            5744: bcd <= 16'h5744;
            5745: bcd <= 16'h5745;
            5746: bcd <= 16'h5746;
            5747: bcd <= 16'h5747;
            5748: bcd <= 16'h5748;
            5749: bcd <= 16'h5749;
            5750: bcd <= 16'h5750;
            5751: bcd <= 16'h5751;
            5752: bcd <= 16'h5752;
            5753: bcd <= 16'h5753;
            5754: bcd <= 16'h5754;
            5755: bcd <= 16'h5755;
            5756: bcd <= 16'h5756;
            5757: bcd <= 16'h5757;
            5758: bcd <= 16'h5758;
            5759: bcd <= 16'h5759;
            5760: bcd <= 16'h5760;
            5761: bcd <= 16'h5761;
            5762: bcd <= 16'h5762;
            5763: bcd <= 16'h5763;
            5764: bcd <= 16'h5764;
            5765: bcd <= 16'h5765;
            5766: bcd <= 16'h5766;
            5767: bcd <= 16'h5767;
            5768: bcd <= 16'h5768;
            5769: bcd <= 16'h5769;
            5770: bcd <= 16'h5770;
            5771: bcd <= 16'h5771;
            5772: bcd <= 16'h5772;
            5773: bcd <= 16'h5773;
            5774: bcd <= 16'h5774;
            5775: bcd <= 16'h5775;
            5776: bcd <= 16'h5776;
            5777: bcd <= 16'h5777;
            5778: bcd <= 16'h5778;
            5779: bcd <= 16'h5779;
            5780: bcd <= 16'h5780;
            5781: bcd <= 16'h5781;
            5782: bcd <= 16'h5782;
            5783: bcd <= 16'h5783;
            5784: bcd <= 16'h5784;
            5785: bcd <= 16'h5785;
            5786: bcd <= 16'h5786;
            5787: bcd <= 16'h5787;
            5788: bcd <= 16'h5788;
            5789: bcd <= 16'h5789;
            5790: bcd <= 16'h5790;
            5791: bcd <= 16'h5791;
            5792: bcd <= 16'h5792;
            5793: bcd <= 16'h5793;
            5794: bcd <= 16'h5794;
            5795: bcd <= 16'h5795;
            5796: bcd <= 16'h5796;
            5797: bcd <= 16'h5797;
            5798: bcd <= 16'h5798;
            5799: bcd <= 16'h5799;
            5800: bcd <= 16'h5800;
            5801: bcd <= 16'h5801;
            5802: bcd <= 16'h5802;
            5803: bcd <= 16'h5803;
            5804: bcd <= 16'h5804;
            5805: bcd <= 16'h5805;
            5806: bcd <= 16'h5806;
            5807: bcd <= 16'h5807;
            5808: bcd <= 16'h5808;
            5809: bcd <= 16'h5809;
            5810: bcd <= 16'h5810;
            5811: bcd <= 16'h5811;
            5812: bcd <= 16'h5812;
            5813: bcd <= 16'h5813;
            5814: bcd <= 16'h5814;
            5815: bcd <= 16'h5815;
            5816: bcd <= 16'h5816;
            5817: bcd <= 16'h5817;
            5818: bcd <= 16'h5818;
            5819: bcd <= 16'h5819;
            5820: bcd <= 16'h5820;
            5821: bcd <= 16'h5821;
            5822: bcd <= 16'h5822;
            5823: bcd <= 16'h5823;
            5824: bcd <= 16'h5824;
            5825: bcd <= 16'h5825;
            5826: bcd <= 16'h5826;
            5827: bcd <= 16'h5827;
            5828: bcd <= 16'h5828;
            5829: bcd <= 16'h5829;
            5830: bcd <= 16'h5830;
            5831: bcd <= 16'h5831;
            5832: bcd <= 16'h5832;
            5833: bcd <= 16'h5833;
            5834: bcd <= 16'h5834;
            5835: bcd <= 16'h5835;
            5836: bcd <= 16'h5836;
            5837: bcd <= 16'h5837;
            5838: bcd <= 16'h5838;
            5839: bcd <= 16'h5839;
            5840: bcd <= 16'h5840;
            5841: bcd <= 16'h5841;
            5842: bcd <= 16'h5842;
            5843: bcd <= 16'h5843;
            5844: bcd <= 16'h5844;
            5845: bcd <= 16'h5845;
            5846: bcd <= 16'h5846;
            5847: bcd <= 16'h5847;
            5848: bcd <= 16'h5848;
            5849: bcd <= 16'h5849;
            5850: bcd <= 16'h5850;
            5851: bcd <= 16'h5851;
            5852: bcd <= 16'h5852;
            5853: bcd <= 16'h5853;
            5854: bcd <= 16'h5854;
            5855: bcd <= 16'h5855;
            5856: bcd <= 16'h5856;
            5857: bcd <= 16'h5857;
            5858: bcd <= 16'h5858;
            5859: bcd <= 16'h5859;
            5860: bcd <= 16'h5860;
            5861: bcd <= 16'h5861;
            5862: bcd <= 16'h5862;
            5863: bcd <= 16'h5863;
            5864: bcd <= 16'h5864;
            5865: bcd <= 16'h5865;
            5866: bcd <= 16'h5866;
            5867: bcd <= 16'h5867;
            5868: bcd <= 16'h5868;
            5869: bcd <= 16'h5869;
            5870: bcd <= 16'h5870;
            5871: bcd <= 16'h5871;
            5872: bcd <= 16'h5872;
            5873: bcd <= 16'h5873;
            5874: bcd <= 16'h5874;
            5875: bcd <= 16'h5875;
            5876: bcd <= 16'h5876;
            5877: bcd <= 16'h5877;
            5878: bcd <= 16'h5878;
            5879: bcd <= 16'h5879;
            5880: bcd <= 16'h5880;
            5881: bcd <= 16'h5881;
            5882: bcd <= 16'h5882;
            5883: bcd <= 16'h5883;
            5884: bcd <= 16'h5884;
            5885: bcd <= 16'h5885;
            5886: bcd <= 16'h5886;
            5887: bcd <= 16'h5887;
            5888: bcd <= 16'h5888;
            5889: bcd <= 16'h5889;
            5890: bcd <= 16'h5890;
            5891: bcd <= 16'h5891;
            5892: bcd <= 16'h5892;
            5893: bcd <= 16'h5893;
            5894: bcd <= 16'h5894;
            5895: bcd <= 16'h5895;
            5896: bcd <= 16'h5896;
            5897: bcd <= 16'h5897;
            5898: bcd <= 16'h5898;
            5899: bcd <= 16'h5899;
            5900: bcd <= 16'h5900;
            5901: bcd <= 16'h5901;
            5902: bcd <= 16'h5902;
            5903: bcd <= 16'h5903;
            5904: bcd <= 16'h5904;
            5905: bcd <= 16'h5905;
            5906: bcd <= 16'h5906;
            5907: bcd <= 16'h5907;
            5908: bcd <= 16'h5908;
            5909: bcd <= 16'h5909;
            5910: bcd <= 16'h5910;
            5911: bcd <= 16'h5911;
            5912: bcd <= 16'h5912;
            5913: bcd <= 16'h5913;
            5914: bcd <= 16'h5914;
            5915: bcd <= 16'h5915;
            5916: bcd <= 16'h5916;
            5917: bcd <= 16'h5917;
            5918: bcd <= 16'h5918;
            5919: bcd <= 16'h5919;
            5920: bcd <= 16'h5920;
            5921: bcd <= 16'h5921;
            5922: bcd <= 16'h5922;
            5923: bcd <= 16'h5923;
            5924: bcd <= 16'h5924;
            5925: bcd <= 16'h5925;
            5926: bcd <= 16'h5926;
            5927: bcd <= 16'h5927;
            5928: bcd <= 16'h5928;
            5929: bcd <= 16'h5929;
            5930: bcd <= 16'h5930;
            5931: bcd <= 16'h5931;
            5932: bcd <= 16'h5932;
            5933: bcd <= 16'h5933;
            5934: bcd <= 16'h5934;
            5935: bcd <= 16'h5935;
            5936: bcd <= 16'h5936;
            5937: bcd <= 16'h5937;
            5938: bcd <= 16'h5938;
            5939: bcd <= 16'h5939;
            5940: bcd <= 16'h5940;
            5941: bcd <= 16'h5941;
            5942: bcd <= 16'h5942;
            5943: bcd <= 16'h5943;
            5944: bcd <= 16'h5944;
            5945: bcd <= 16'h5945;
            5946: bcd <= 16'h5946;
            5947: bcd <= 16'h5947;
            5948: bcd <= 16'h5948;
            5949: bcd <= 16'h5949;
            5950: bcd <= 16'h5950;
            5951: bcd <= 16'h5951;
            5952: bcd <= 16'h5952;
            5953: bcd <= 16'h5953;
            5954: bcd <= 16'h5954;
            5955: bcd <= 16'h5955;
            5956: bcd <= 16'h5956;
            5957: bcd <= 16'h5957;
            5958: bcd <= 16'h5958;
            5959: bcd <= 16'h5959;
            5960: bcd <= 16'h5960;
            5961: bcd <= 16'h5961;
            5962: bcd <= 16'h5962;
            5963: bcd <= 16'h5963;
            5964: bcd <= 16'h5964;
            5965: bcd <= 16'h5965;
            5966: bcd <= 16'h5966;
            5967: bcd <= 16'h5967;
            5968: bcd <= 16'h5968;
            5969: bcd <= 16'h5969;
            5970: bcd <= 16'h5970;
            5971: bcd <= 16'h5971;
            5972: bcd <= 16'h5972;
            5973: bcd <= 16'h5973;
            5974: bcd <= 16'h5974;
            5975: bcd <= 16'h5975;
            5976: bcd <= 16'h5976;
            5977: bcd <= 16'h5977;
            5978: bcd <= 16'h5978;
            5979: bcd <= 16'h5979;
            5980: bcd <= 16'h5980;
            5981: bcd <= 16'h5981;
            5982: bcd <= 16'h5982;
            5983: bcd <= 16'h5983;
            5984: bcd <= 16'h5984;
            5985: bcd <= 16'h5985;
            5986: bcd <= 16'h5986;
            5987: bcd <= 16'h5987;
            5988: bcd <= 16'h5988;
            5989: bcd <= 16'h5989;
            5990: bcd <= 16'h5990;
            5991: bcd <= 16'h5991;
            5992: bcd <= 16'h5992;
            5993: bcd <= 16'h5993;
            5994: bcd <= 16'h5994;
            5995: bcd <= 16'h5995;
            5996: bcd <= 16'h5996;
            5997: bcd <= 16'h5997;
            5998: bcd <= 16'h5998;
            5999: bcd <= 16'h5999;
            6000: bcd <= 16'h6000;
            6001: bcd <= 16'h6001;
            6002: bcd <= 16'h6002;
            6003: bcd <= 16'h6003;
            6004: bcd <= 16'h6004;
            6005: bcd <= 16'h6005;
            6006: bcd <= 16'h6006;
            6007: bcd <= 16'h6007;
            6008: bcd <= 16'h6008;
            6009: bcd <= 16'h6009;
            6010: bcd <= 16'h6010;
            6011: bcd <= 16'h6011;
            6012: bcd <= 16'h6012;
            6013: bcd <= 16'h6013;
            6014: bcd <= 16'h6014;
            6015: bcd <= 16'h6015;
            6016: bcd <= 16'h6016;
            6017: bcd <= 16'h6017;
            6018: bcd <= 16'h6018;
            6019: bcd <= 16'h6019;
            6020: bcd <= 16'h6020;
            6021: bcd <= 16'h6021;
            6022: bcd <= 16'h6022;
            6023: bcd <= 16'h6023;
            6024: bcd <= 16'h6024;
            6025: bcd <= 16'h6025;
            6026: bcd <= 16'h6026;
            6027: bcd <= 16'h6027;
            6028: bcd <= 16'h6028;
            6029: bcd <= 16'h6029;
            6030: bcd <= 16'h6030;
            6031: bcd <= 16'h6031;
            6032: bcd <= 16'h6032;
            6033: bcd <= 16'h6033;
            6034: bcd <= 16'h6034;
            6035: bcd <= 16'h6035;
            6036: bcd <= 16'h6036;
            6037: bcd <= 16'h6037;
            6038: bcd <= 16'h6038;
            6039: bcd <= 16'h6039;
            6040: bcd <= 16'h6040;
            6041: bcd <= 16'h6041;
            6042: bcd <= 16'h6042;
            6043: bcd <= 16'h6043;
            6044: bcd <= 16'h6044;
            6045: bcd <= 16'h6045;
            6046: bcd <= 16'h6046;
            6047: bcd <= 16'h6047;
            6048: bcd <= 16'h6048;
            6049: bcd <= 16'h6049;
            6050: bcd <= 16'h6050;
            6051: bcd <= 16'h6051;
            6052: bcd <= 16'h6052;
            6053: bcd <= 16'h6053;
            6054: bcd <= 16'h6054;
            6055: bcd <= 16'h6055;
            6056: bcd <= 16'h6056;
            6057: bcd <= 16'h6057;
            6058: bcd <= 16'h6058;
            6059: bcd <= 16'h6059;
            6060: bcd <= 16'h6060;
            6061: bcd <= 16'h6061;
            6062: bcd <= 16'h6062;
            6063: bcd <= 16'h6063;
            6064: bcd <= 16'h6064;
            6065: bcd <= 16'h6065;
            6066: bcd <= 16'h6066;
            6067: bcd <= 16'h6067;
            6068: bcd <= 16'h6068;
            6069: bcd <= 16'h6069;
            6070: bcd <= 16'h6070;
            6071: bcd <= 16'h6071;
            6072: bcd <= 16'h6072;
            6073: bcd <= 16'h6073;
            6074: bcd <= 16'h6074;
            6075: bcd <= 16'h6075;
            6076: bcd <= 16'h6076;
            6077: bcd <= 16'h6077;
            6078: bcd <= 16'h6078;
            6079: bcd <= 16'h6079;
            6080: bcd <= 16'h6080;
            6081: bcd <= 16'h6081;
            6082: bcd <= 16'h6082;
            6083: bcd <= 16'h6083;
            6084: bcd <= 16'h6084;
            6085: bcd <= 16'h6085;
            6086: bcd <= 16'h6086;
            6087: bcd <= 16'h6087;
            6088: bcd <= 16'h6088;
            6089: bcd <= 16'h6089;
            6090: bcd <= 16'h6090;
            6091: bcd <= 16'h6091;
            6092: bcd <= 16'h6092;
            6093: bcd <= 16'h6093;
            6094: bcd <= 16'h6094;
            6095: bcd <= 16'h6095;
            6096: bcd <= 16'h6096;
            6097: bcd <= 16'h6097;
            6098: bcd <= 16'h6098;
            6099: bcd <= 16'h6099;
            6100: bcd <= 16'h6100;
            6101: bcd <= 16'h6101;
            6102: bcd <= 16'h6102;
            6103: bcd <= 16'h6103;
            6104: bcd <= 16'h6104;
            6105: bcd <= 16'h6105;
            6106: bcd <= 16'h6106;
            6107: bcd <= 16'h6107;
            6108: bcd <= 16'h6108;
            6109: bcd <= 16'h6109;
            6110: bcd <= 16'h6110;
            6111: bcd <= 16'h6111;
            6112: bcd <= 16'h6112;
            6113: bcd <= 16'h6113;
            6114: bcd <= 16'h6114;
            6115: bcd <= 16'h6115;
            6116: bcd <= 16'h6116;
            6117: bcd <= 16'h6117;
            6118: bcd <= 16'h6118;
            6119: bcd <= 16'h6119;
            6120: bcd <= 16'h6120;
            6121: bcd <= 16'h6121;
            6122: bcd <= 16'h6122;
            6123: bcd <= 16'h6123;
            6124: bcd <= 16'h6124;
            6125: bcd <= 16'h6125;
            6126: bcd <= 16'h6126;
            6127: bcd <= 16'h6127;
            6128: bcd <= 16'h6128;
            6129: bcd <= 16'h6129;
            6130: bcd <= 16'h6130;
            6131: bcd <= 16'h6131;
            6132: bcd <= 16'h6132;
            6133: bcd <= 16'h6133;
            6134: bcd <= 16'h6134;
            6135: bcd <= 16'h6135;
            6136: bcd <= 16'h6136;
            6137: bcd <= 16'h6137;
            6138: bcd <= 16'h6138;
            6139: bcd <= 16'h6139;
            6140: bcd <= 16'h6140;
            6141: bcd <= 16'h6141;
            6142: bcd <= 16'h6142;
            6143: bcd <= 16'h6143;
            6144: bcd <= 16'h6144;
            6145: bcd <= 16'h6145;
            6146: bcd <= 16'h6146;
            6147: bcd <= 16'h6147;
            6148: bcd <= 16'h6148;
            6149: bcd <= 16'h6149;
            6150: bcd <= 16'h6150;
            6151: bcd <= 16'h6151;
            6152: bcd <= 16'h6152;
            6153: bcd <= 16'h6153;
            6154: bcd <= 16'h6154;
            6155: bcd <= 16'h6155;
            6156: bcd <= 16'h6156;
            6157: bcd <= 16'h6157;
            6158: bcd <= 16'h6158;
            6159: bcd <= 16'h6159;
            6160: bcd <= 16'h6160;
            6161: bcd <= 16'h6161;
            6162: bcd <= 16'h6162;
            6163: bcd <= 16'h6163;
            6164: bcd <= 16'h6164;
            6165: bcd <= 16'h6165;
            6166: bcd <= 16'h6166;
            6167: bcd <= 16'h6167;
            6168: bcd <= 16'h6168;
            6169: bcd <= 16'h6169;
            6170: bcd <= 16'h6170;
            6171: bcd <= 16'h6171;
            6172: bcd <= 16'h6172;
            6173: bcd <= 16'h6173;
            6174: bcd <= 16'h6174;
            6175: bcd <= 16'h6175;
            6176: bcd <= 16'h6176;
            6177: bcd <= 16'h6177;
            6178: bcd <= 16'h6178;
            6179: bcd <= 16'h6179;
            6180: bcd <= 16'h6180;
            6181: bcd <= 16'h6181;
            6182: bcd <= 16'h6182;
            6183: bcd <= 16'h6183;
            6184: bcd <= 16'h6184;
            6185: bcd <= 16'h6185;
            6186: bcd <= 16'h6186;
            6187: bcd <= 16'h6187;
            6188: bcd <= 16'h6188;
            6189: bcd <= 16'h6189;
            6190: bcd <= 16'h6190;
            6191: bcd <= 16'h6191;
            6192: bcd <= 16'h6192;
            6193: bcd <= 16'h6193;
            6194: bcd <= 16'h6194;
            6195: bcd <= 16'h6195;
            6196: bcd <= 16'h6196;
            6197: bcd <= 16'h6197;
            6198: bcd <= 16'h6198;
            6199: bcd <= 16'h6199;
            6200: bcd <= 16'h6200;
            6201: bcd <= 16'h6201;
            6202: bcd <= 16'h6202;
            6203: bcd <= 16'h6203;
            6204: bcd <= 16'h6204;
            6205: bcd <= 16'h6205;
            6206: bcd <= 16'h6206;
            6207: bcd <= 16'h6207;
            6208: bcd <= 16'h6208;
            6209: bcd <= 16'h6209;
            6210: bcd <= 16'h6210;
            6211: bcd <= 16'h6211;
            6212: bcd <= 16'h6212;
            6213: bcd <= 16'h6213;
            6214: bcd <= 16'h6214;
            6215: bcd <= 16'h6215;
            6216: bcd <= 16'h6216;
            6217: bcd <= 16'h6217;
            6218: bcd <= 16'h6218;
            6219: bcd <= 16'h6219;
            6220: bcd <= 16'h6220;
            6221: bcd <= 16'h6221;
            6222: bcd <= 16'h6222;
            6223: bcd <= 16'h6223;
            6224: bcd <= 16'h6224;
            6225: bcd <= 16'h6225;
            6226: bcd <= 16'h6226;
            6227: bcd <= 16'h6227;
            6228: bcd <= 16'h6228;
            6229: bcd <= 16'h6229;
            6230: bcd <= 16'h6230;
            6231: bcd <= 16'h6231;
            6232: bcd <= 16'h6232;
            6233: bcd <= 16'h6233;
            6234: bcd <= 16'h6234;
            6235: bcd <= 16'h6235;
            6236: bcd <= 16'h6236;
            6237: bcd <= 16'h6237;
            6238: bcd <= 16'h6238;
            6239: bcd <= 16'h6239;
            6240: bcd <= 16'h6240;
            6241: bcd <= 16'h6241;
            6242: bcd <= 16'h6242;
            6243: bcd <= 16'h6243;
            6244: bcd <= 16'h6244;
            6245: bcd <= 16'h6245;
            6246: bcd <= 16'h6246;
            6247: bcd <= 16'h6247;
            6248: bcd <= 16'h6248;
            6249: bcd <= 16'h6249;
            6250: bcd <= 16'h6250;
            6251: bcd <= 16'h6251;
            6252: bcd <= 16'h6252;
            6253: bcd <= 16'h6253;
            6254: bcd <= 16'h6254;
            6255: bcd <= 16'h6255;
            6256: bcd <= 16'h6256;
            6257: bcd <= 16'h6257;
            6258: bcd <= 16'h6258;
            6259: bcd <= 16'h6259;
            6260: bcd <= 16'h6260;
            6261: bcd <= 16'h6261;
            6262: bcd <= 16'h6262;
            6263: bcd <= 16'h6263;
            6264: bcd <= 16'h6264;
            6265: bcd <= 16'h6265;
            6266: bcd <= 16'h6266;
            6267: bcd <= 16'h6267;
            6268: bcd <= 16'h6268;
            6269: bcd <= 16'h6269;
            6270: bcd <= 16'h6270;
            6271: bcd <= 16'h6271;
            6272: bcd <= 16'h6272;
            6273: bcd <= 16'h6273;
            6274: bcd <= 16'h6274;
            6275: bcd <= 16'h6275;
            6276: bcd <= 16'h6276;
            6277: bcd <= 16'h6277;
            6278: bcd <= 16'h6278;
            6279: bcd <= 16'h6279;
            6280: bcd <= 16'h6280;
            6281: bcd <= 16'h6281;
            6282: bcd <= 16'h6282;
            6283: bcd <= 16'h6283;
            6284: bcd <= 16'h6284;
            6285: bcd <= 16'h6285;
            6286: bcd <= 16'h6286;
            6287: bcd <= 16'h6287;
            6288: bcd <= 16'h6288;
            6289: bcd <= 16'h6289;
            6290: bcd <= 16'h6290;
            6291: bcd <= 16'h6291;
            6292: bcd <= 16'h6292;
            6293: bcd <= 16'h6293;
            6294: bcd <= 16'h6294;
            6295: bcd <= 16'h6295;
            6296: bcd <= 16'h6296;
            6297: bcd <= 16'h6297;
            6298: bcd <= 16'h6298;
            6299: bcd <= 16'h6299;
            6300: bcd <= 16'h6300;
            6301: bcd <= 16'h6301;
            6302: bcd <= 16'h6302;
            6303: bcd <= 16'h6303;
            6304: bcd <= 16'h6304;
            6305: bcd <= 16'h6305;
            6306: bcd <= 16'h6306;
            6307: bcd <= 16'h6307;
            6308: bcd <= 16'h6308;
            6309: bcd <= 16'h6309;
            6310: bcd <= 16'h6310;
            6311: bcd <= 16'h6311;
            6312: bcd <= 16'h6312;
            6313: bcd <= 16'h6313;
            6314: bcd <= 16'h6314;
            6315: bcd <= 16'h6315;
            6316: bcd <= 16'h6316;
            6317: bcd <= 16'h6317;
            6318: bcd <= 16'h6318;
            6319: bcd <= 16'h6319;
            6320: bcd <= 16'h6320;
            6321: bcd <= 16'h6321;
            6322: bcd <= 16'h6322;
            6323: bcd <= 16'h6323;
            6324: bcd <= 16'h6324;
            6325: bcd <= 16'h6325;
            6326: bcd <= 16'h6326;
            6327: bcd <= 16'h6327;
            6328: bcd <= 16'h6328;
            6329: bcd <= 16'h6329;
            6330: bcd <= 16'h6330;
            6331: bcd <= 16'h6331;
            6332: bcd <= 16'h6332;
            6333: bcd <= 16'h6333;
            6334: bcd <= 16'h6334;
            6335: bcd <= 16'h6335;
            6336: bcd <= 16'h6336;
            6337: bcd <= 16'h6337;
            6338: bcd <= 16'h6338;
            6339: bcd <= 16'h6339;
            6340: bcd <= 16'h6340;
            6341: bcd <= 16'h6341;
            6342: bcd <= 16'h6342;
            6343: bcd <= 16'h6343;
            6344: bcd <= 16'h6344;
            6345: bcd <= 16'h6345;
            6346: bcd <= 16'h6346;
            6347: bcd <= 16'h6347;
            6348: bcd <= 16'h6348;
            6349: bcd <= 16'h6349;
            6350: bcd <= 16'h6350;
            6351: bcd <= 16'h6351;
            6352: bcd <= 16'h6352;
            6353: bcd <= 16'h6353;
            6354: bcd <= 16'h6354;
            6355: bcd <= 16'h6355;
            6356: bcd <= 16'h6356;
            6357: bcd <= 16'h6357;
            6358: bcd <= 16'h6358;
            6359: bcd <= 16'h6359;
            6360: bcd <= 16'h6360;
            6361: bcd <= 16'h6361;
            6362: bcd <= 16'h6362;
            6363: bcd <= 16'h6363;
            6364: bcd <= 16'h6364;
            6365: bcd <= 16'h6365;
            6366: bcd <= 16'h6366;
            6367: bcd <= 16'h6367;
            6368: bcd <= 16'h6368;
            6369: bcd <= 16'h6369;
            6370: bcd <= 16'h6370;
            6371: bcd <= 16'h6371;
            6372: bcd <= 16'h6372;
            6373: bcd <= 16'h6373;
            6374: bcd <= 16'h6374;
            6375: bcd <= 16'h6375;
            6376: bcd <= 16'h6376;
            6377: bcd <= 16'h6377;
            6378: bcd <= 16'h6378;
            6379: bcd <= 16'h6379;
            6380: bcd <= 16'h6380;
            6381: bcd <= 16'h6381;
            6382: bcd <= 16'h6382;
            6383: bcd <= 16'h6383;
            6384: bcd <= 16'h6384;
            6385: bcd <= 16'h6385;
            6386: bcd <= 16'h6386;
            6387: bcd <= 16'h6387;
            6388: bcd <= 16'h6388;
            6389: bcd <= 16'h6389;
            6390: bcd <= 16'h6390;
            6391: bcd <= 16'h6391;
            6392: bcd <= 16'h6392;
            6393: bcd <= 16'h6393;
            6394: bcd <= 16'h6394;
            6395: bcd <= 16'h6395;
            6396: bcd <= 16'h6396;
            6397: bcd <= 16'h6397;
            6398: bcd <= 16'h6398;
            6399: bcd <= 16'h6399;
            6400: bcd <= 16'h6400;
            6401: bcd <= 16'h6401;
            6402: bcd <= 16'h6402;
            6403: bcd <= 16'h6403;
            6404: bcd <= 16'h6404;
            6405: bcd <= 16'h6405;
            6406: bcd <= 16'h6406;
            6407: bcd <= 16'h6407;
            6408: bcd <= 16'h6408;
            6409: bcd <= 16'h6409;
            6410: bcd <= 16'h6410;
            6411: bcd <= 16'h6411;
            6412: bcd <= 16'h6412;
            6413: bcd <= 16'h6413;
            6414: bcd <= 16'h6414;
            6415: bcd <= 16'h6415;
            6416: bcd <= 16'h6416;
            6417: bcd <= 16'h6417;
            6418: bcd <= 16'h6418;
            6419: bcd <= 16'h6419;
            6420: bcd <= 16'h6420;
            6421: bcd <= 16'h6421;
            6422: bcd <= 16'h6422;
            6423: bcd <= 16'h6423;
            6424: bcd <= 16'h6424;
            6425: bcd <= 16'h6425;
            6426: bcd <= 16'h6426;
            6427: bcd <= 16'h6427;
            6428: bcd <= 16'h6428;
            6429: bcd <= 16'h6429;
            6430: bcd <= 16'h6430;
            6431: bcd <= 16'h6431;
            6432: bcd <= 16'h6432;
            6433: bcd <= 16'h6433;
            6434: bcd <= 16'h6434;
            6435: bcd <= 16'h6435;
            6436: bcd <= 16'h6436;
            6437: bcd <= 16'h6437;
            6438: bcd <= 16'h6438;
            6439: bcd <= 16'h6439;
            6440: bcd <= 16'h6440;
            6441: bcd <= 16'h6441;
            6442: bcd <= 16'h6442;
            6443: bcd <= 16'h6443;
            6444: bcd <= 16'h6444;
            6445: bcd <= 16'h6445;
            6446: bcd <= 16'h6446;
            6447: bcd <= 16'h6447;
            6448: bcd <= 16'h6448;
            6449: bcd <= 16'h6449;
            6450: bcd <= 16'h6450;
            6451: bcd <= 16'h6451;
            6452: bcd <= 16'h6452;
            6453: bcd <= 16'h6453;
            6454: bcd <= 16'h6454;
            6455: bcd <= 16'h6455;
            6456: bcd <= 16'h6456;
            6457: bcd <= 16'h6457;
            6458: bcd <= 16'h6458;
            6459: bcd <= 16'h6459;
            6460: bcd <= 16'h6460;
            6461: bcd <= 16'h6461;
            6462: bcd <= 16'h6462;
            6463: bcd <= 16'h6463;
            6464: bcd <= 16'h6464;
            6465: bcd <= 16'h6465;
            6466: bcd <= 16'h6466;
            6467: bcd <= 16'h6467;
            6468: bcd <= 16'h6468;
            6469: bcd <= 16'h6469;
            6470: bcd <= 16'h6470;
            6471: bcd <= 16'h6471;
            6472: bcd <= 16'h6472;
            6473: bcd <= 16'h6473;
            6474: bcd <= 16'h6474;
            6475: bcd <= 16'h6475;
            6476: bcd <= 16'h6476;
            6477: bcd <= 16'h6477;
            6478: bcd <= 16'h6478;
            6479: bcd <= 16'h6479;
            6480: bcd <= 16'h6480;
            6481: bcd <= 16'h6481;
            6482: bcd <= 16'h6482;
            6483: bcd <= 16'h6483;
            6484: bcd <= 16'h6484;
            6485: bcd <= 16'h6485;
            6486: bcd <= 16'h6486;
            6487: bcd <= 16'h6487;
            6488: bcd <= 16'h6488;
            6489: bcd <= 16'h6489;
            6490: bcd <= 16'h6490;
            6491: bcd <= 16'h6491;
            6492: bcd <= 16'h6492;
            6493: bcd <= 16'h6493;
            6494: bcd <= 16'h6494;
            6495: bcd <= 16'h6495;
            6496: bcd <= 16'h6496;
            6497: bcd <= 16'h6497;
            6498: bcd <= 16'h6498;
            6499: bcd <= 16'h6499;
            6500: bcd <= 16'h6500;
            6501: bcd <= 16'h6501;
            6502: bcd <= 16'h6502;
            6503: bcd <= 16'h6503;
            6504: bcd <= 16'h6504;
            6505: bcd <= 16'h6505;
            6506: bcd <= 16'h6506;
            6507: bcd <= 16'h6507;
            6508: bcd <= 16'h6508;
            6509: bcd <= 16'h6509;
            6510: bcd <= 16'h6510;
            6511: bcd <= 16'h6511;
            6512: bcd <= 16'h6512;
            6513: bcd <= 16'h6513;
            6514: bcd <= 16'h6514;
            6515: bcd <= 16'h6515;
            6516: bcd <= 16'h6516;
            6517: bcd <= 16'h6517;
            6518: bcd <= 16'h6518;
            6519: bcd <= 16'h6519;
            6520: bcd <= 16'h6520;
            6521: bcd <= 16'h6521;
            6522: bcd <= 16'h6522;
            6523: bcd <= 16'h6523;
            6524: bcd <= 16'h6524;
            6525: bcd <= 16'h6525;
            6526: bcd <= 16'h6526;
            6527: bcd <= 16'h6527;
            6528: bcd <= 16'h6528;
            6529: bcd <= 16'h6529;
            6530: bcd <= 16'h6530;
            6531: bcd <= 16'h6531;
            6532: bcd <= 16'h6532;
            6533: bcd <= 16'h6533;
            6534: bcd <= 16'h6534;
            6535: bcd <= 16'h6535;
            6536: bcd <= 16'h6536;
            6537: bcd <= 16'h6537;
            6538: bcd <= 16'h6538;
            6539: bcd <= 16'h6539;
            6540: bcd <= 16'h6540;
            6541: bcd <= 16'h6541;
            6542: bcd <= 16'h6542;
            6543: bcd <= 16'h6543;
            6544: bcd <= 16'h6544;
            6545: bcd <= 16'h6545;
            6546: bcd <= 16'h6546;
            6547: bcd <= 16'h6547;
            6548: bcd <= 16'h6548;
            6549: bcd <= 16'h6549;
            6550: bcd <= 16'h6550;
            6551: bcd <= 16'h6551;
            6552: bcd <= 16'h6552;
            6553: bcd <= 16'h6553;
            6554: bcd <= 16'h6554;
            6555: bcd <= 16'h6555;
            6556: bcd <= 16'h6556;
            6557: bcd <= 16'h6557;
            6558: bcd <= 16'h6558;
            6559: bcd <= 16'h6559;
            6560: bcd <= 16'h6560;
            6561: bcd <= 16'h6561;
            6562: bcd <= 16'h6562;
            6563: bcd <= 16'h6563;
            6564: bcd <= 16'h6564;
            6565: bcd <= 16'h6565;
            6566: bcd <= 16'h6566;
            6567: bcd <= 16'h6567;
            6568: bcd <= 16'h6568;
            6569: bcd <= 16'h6569;
            6570: bcd <= 16'h6570;
            6571: bcd <= 16'h6571;
            6572: bcd <= 16'h6572;
            6573: bcd <= 16'h6573;
            6574: bcd <= 16'h6574;
            6575: bcd <= 16'h6575;
            6576: bcd <= 16'h6576;
            6577: bcd <= 16'h6577;
            6578: bcd <= 16'h6578;
            6579: bcd <= 16'h6579;
            6580: bcd <= 16'h6580;
            6581: bcd <= 16'h6581;
            6582: bcd <= 16'h6582;
            6583: bcd <= 16'h6583;
            6584: bcd <= 16'h6584;
            6585: bcd <= 16'h6585;
            6586: bcd <= 16'h6586;
            6587: bcd <= 16'h6587;
            6588: bcd <= 16'h6588;
            6589: bcd <= 16'h6589;
            6590: bcd <= 16'h6590;
            6591: bcd <= 16'h6591;
            6592: bcd <= 16'h6592;
            6593: bcd <= 16'h6593;
            6594: bcd <= 16'h6594;
            6595: bcd <= 16'h6595;
            6596: bcd <= 16'h6596;
            6597: bcd <= 16'h6597;
            6598: bcd <= 16'h6598;
            6599: bcd <= 16'h6599;
            6600: bcd <= 16'h6600;
            6601: bcd <= 16'h6601;
            6602: bcd <= 16'h6602;
            6603: bcd <= 16'h6603;
            6604: bcd <= 16'h6604;
            6605: bcd <= 16'h6605;
            6606: bcd <= 16'h6606;
            6607: bcd <= 16'h6607;
            6608: bcd <= 16'h6608;
            6609: bcd <= 16'h6609;
            6610: bcd <= 16'h6610;
            6611: bcd <= 16'h6611;
            6612: bcd <= 16'h6612;
            6613: bcd <= 16'h6613;
            6614: bcd <= 16'h6614;
            6615: bcd <= 16'h6615;
            6616: bcd <= 16'h6616;
            6617: bcd <= 16'h6617;
            6618: bcd <= 16'h6618;
            6619: bcd <= 16'h6619;
            6620: bcd <= 16'h6620;
            6621: bcd <= 16'h6621;
            6622: bcd <= 16'h6622;
            6623: bcd <= 16'h6623;
            6624: bcd <= 16'h6624;
            6625: bcd <= 16'h6625;
            6626: bcd <= 16'h6626;
            6627: bcd <= 16'h6627;
            6628: bcd <= 16'h6628;
            6629: bcd <= 16'h6629;
            6630: bcd <= 16'h6630;
            6631: bcd <= 16'h6631;
            6632: bcd <= 16'h6632;
            6633: bcd <= 16'h6633;
            6634: bcd <= 16'h6634;
            6635: bcd <= 16'h6635;
            6636: bcd <= 16'h6636;
            6637: bcd <= 16'h6637;
            6638: bcd <= 16'h6638;
            6639: bcd <= 16'h6639;
            6640: bcd <= 16'h6640;
            6641: bcd <= 16'h6641;
            6642: bcd <= 16'h6642;
            6643: bcd <= 16'h6643;
            6644: bcd <= 16'h6644;
            6645: bcd <= 16'h6645;
            6646: bcd <= 16'h6646;
            6647: bcd <= 16'h6647;
            6648: bcd <= 16'h6648;
            6649: bcd <= 16'h6649;
            6650: bcd <= 16'h6650;
            6651: bcd <= 16'h6651;
            6652: bcd <= 16'h6652;
            6653: bcd <= 16'h6653;
            6654: bcd <= 16'h6654;
            6655: bcd <= 16'h6655;
            6656: bcd <= 16'h6656;
            6657: bcd <= 16'h6657;
            6658: bcd <= 16'h6658;
            6659: bcd <= 16'h6659;
            6660: bcd <= 16'h6660;
            6661: bcd <= 16'h6661;
            6662: bcd <= 16'h6662;
            6663: bcd <= 16'h6663;
            6664: bcd <= 16'h6664;
            6665: bcd <= 16'h6665;
            6666: bcd <= 16'h6666;
            6667: bcd <= 16'h6667;
            6668: bcd <= 16'h6668;
            6669: bcd <= 16'h6669;
            6670: bcd <= 16'h6670;
            6671: bcd <= 16'h6671;
            6672: bcd <= 16'h6672;
            6673: bcd <= 16'h6673;
            6674: bcd <= 16'h6674;
            6675: bcd <= 16'h6675;
            6676: bcd <= 16'h6676;
            6677: bcd <= 16'h6677;
            6678: bcd <= 16'h6678;
            6679: bcd <= 16'h6679;
            6680: bcd <= 16'h6680;
            6681: bcd <= 16'h6681;
            6682: bcd <= 16'h6682;
            6683: bcd <= 16'h6683;
            6684: bcd <= 16'h6684;
            6685: bcd <= 16'h6685;
            6686: bcd <= 16'h6686;
            6687: bcd <= 16'h6687;
            6688: bcd <= 16'h6688;
            6689: bcd <= 16'h6689;
            6690: bcd <= 16'h6690;
            6691: bcd <= 16'h6691;
            6692: bcd <= 16'h6692;
            6693: bcd <= 16'h6693;
            6694: bcd <= 16'h6694;
            6695: bcd <= 16'h6695;
            6696: bcd <= 16'h6696;
            6697: bcd <= 16'h6697;
            6698: bcd <= 16'h6698;
            6699: bcd <= 16'h6699;
            6700: bcd <= 16'h6700;
            6701: bcd <= 16'h6701;
            6702: bcd <= 16'h6702;
            6703: bcd <= 16'h6703;
            6704: bcd <= 16'h6704;
            6705: bcd <= 16'h6705;
            6706: bcd <= 16'h6706;
            6707: bcd <= 16'h6707;
            6708: bcd <= 16'h6708;
            6709: bcd <= 16'h6709;
            6710: bcd <= 16'h6710;
            6711: bcd <= 16'h6711;
            6712: bcd <= 16'h6712;
            6713: bcd <= 16'h6713;
            6714: bcd <= 16'h6714;
            6715: bcd <= 16'h6715;
            6716: bcd <= 16'h6716;
            6717: bcd <= 16'h6717;
            6718: bcd <= 16'h6718;
            6719: bcd <= 16'h6719;
            6720: bcd <= 16'h6720;
            6721: bcd <= 16'h6721;
            6722: bcd <= 16'h6722;
            6723: bcd <= 16'h6723;
            6724: bcd <= 16'h6724;
            6725: bcd <= 16'h6725;
            6726: bcd <= 16'h6726;
            6727: bcd <= 16'h6727;
            6728: bcd <= 16'h6728;
            6729: bcd <= 16'h6729;
            6730: bcd <= 16'h6730;
            6731: bcd <= 16'h6731;
            6732: bcd <= 16'h6732;
            6733: bcd <= 16'h6733;
            6734: bcd <= 16'h6734;
            6735: bcd <= 16'h6735;
            6736: bcd <= 16'h6736;
            6737: bcd <= 16'h6737;
            6738: bcd <= 16'h6738;
            6739: bcd <= 16'h6739;
            6740: bcd <= 16'h6740;
            6741: bcd <= 16'h6741;
            6742: bcd <= 16'h6742;
            6743: bcd <= 16'h6743;
            6744: bcd <= 16'h6744;
            6745: bcd <= 16'h6745;
            6746: bcd <= 16'h6746;
            6747: bcd <= 16'h6747;
            6748: bcd <= 16'h6748;
            6749: bcd <= 16'h6749;
            6750: bcd <= 16'h6750;
            6751: bcd <= 16'h6751;
            6752: bcd <= 16'h6752;
            6753: bcd <= 16'h6753;
            6754: bcd <= 16'h6754;
            6755: bcd <= 16'h6755;
            6756: bcd <= 16'h6756;
            6757: bcd <= 16'h6757;
            6758: bcd <= 16'h6758;
            6759: bcd <= 16'h6759;
            6760: bcd <= 16'h6760;
            6761: bcd <= 16'h6761;
            6762: bcd <= 16'h6762;
            6763: bcd <= 16'h6763;
            6764: bcd <= 16'h6764;
            6765: bcd <= 16'h6765;
            6766: bcd <= 16'h6766;
            6767: bcd <= 16'h6767;
            6768: bcd <= 16'h6768;
            6769: bcd <= 16'h6769;
            6770: bcd <= 16'h6770;
            6771: bcd <= 16'h6771;
            6772: bcd <= 16'h6772;
            6773: bcd <= 16'h6773;
            6774: bcd <= 16'h6774;
            6775: bcd <= 16'h6775;
            6776: bcd <= 16'h6776;
            6777: bcd <= 16'h6777;
            6778: bcd <= 16'h6778;
            6779: bcd <= 16'h6779;
            6780: bcd <= 16'h6780;
            6781: bcd <= 16'h6781;
            6782: bcd <= 16'h6782;
            6783: bcd <= 16'h6783;
            6784: bcd <= 16'h6784;
            6785: bcd <= 16'h6785;
            6786: bcd <= 16'h6786;
            6787: bcd <= 16'h6787;
            6788: bcd <= 16'h6788;
            6789: bcd <= 16'h6789;
            6790: bcd <= 16'h6790;
            6791: bcd <= 16'h6791;
            6792: bcd <= 16'h6792;
            6793: bcd <= 16'h6793;
            6794: bcd <= 16'h6794;
            6795: bcd <= 16'h6795;
            6796: bcd <= 16'h6796;
            6797: bcd <= 16'h6797;
            6798: bcd <= 16'h6798;
            6799: bcd <= 16'h6799;
            6800: bcd <= 16'h6800;
            6801: bcd <= 16'h6801;
            6802: bcd <= 16'h6802;
            6803: bcd <= 16'h6803;
            6804: bcd <= 16'h6804;
            6805: bcd <= 16'h6805;
            6806: bcd <= 16'h6806;
            6807: bcd <= 16'h6807;
            6808: bcd <= 16'h6808;
            6809: bcd <= 16'h6809;
            6810: bcd <= 16'h6810;
            6811: bcd <= 16'h6811;
            6812: bcd <= 16'h6812;
            6813: bcd <= 16'h6813;
            6814: bcd <= 16'h6814;
            6815: bcd <= 16'h6815;
            6816: bcd <= 16'h6816;
            6817: bcd <= 16'h6817;
            6818: bcd <= 16'h6818;
            6819: bcd <= 16'h6819;
            6820: bcd <= 16'h6820;
            6821: bcd <= 16'h6821;
            6822: bcd <= 16'h6822;
            6823: bcd <= 16'h6823;
            6824: bcd <= 16'h6824;
            6825: bcd <= 16'h6825;
            6826: bcd <= 16'h6826;
            6827: bcd <= 16'h6827;
            6828: bcd <= 16'h6828;
            6829: bcd <= 16'h6829;
            6830: bcd <= 16'h6830;
            6831: bcd <= 16'h6831;
            6832: bcd <= 16'h6832;
            6833: bcd <= 16'h6833;
            6834: bcd <= 16'h6834;
            6835: bcd <= 16'h6835;
            6836: bcd <= 16'h6836;
            6837: bcd <= 16'h6837;
            6838: bcd <= 16'h6838;
            6839: bcd <= 16'h6839;
            6840: bcd <= 16'h6840;
            6841: bcd <= 16'h6841;
            6842: bcd <= 16'h6842;
            6843: bcd <= 16'h6843;
            6844: bcd <= 16'h6844;
            6845: bcd <= 16'h6845;
            6846: bcd <= 16'h6846;
            6847: bcd <= 16'h6847;
            6848: bcd <= 16'h6848;
            6849: bcd <= 16'h6849;
            6850: bcd <= 16'h6850;
            6851: bcd <= 16'h6851;
            6852: bcd <= 16'h6852;
            6853: bcd <= 16'h6853;
            6854: bcd <= 16'h6854;
            6855: bcd <= 16'h6855;
            6856: bcd <= 16'h6856;
            6857: bcd <= 16'h6857;
            6858: bcd <= 16'h6858;
            6859: bcd <= 16'h6859;
            6860: bcd <= 16'h6860;
            6861: bcd <= 16'h6861;
            6862: bcd <= 16'h6862;
            6863: bcd <= 16'h6863;
            6864: bcd <= 16'h6864;
            6865: bcd <= 16'h6865;
            6866: bcd <= 16'h6866;
            6867: bcd <= 16'h6867;
            6868: bcd <= 16'h6868;
            6869: bcd <= 16'h6869;
            6870: bcd <= 16'h6870;
            6871: bcd <= 16'h6871;
            6872: bcd <= 16'h6872;
            6873: bcd <= 16'h6873;
            6874: bcd <= 16'h6874;
            6875: bcd <= 16'h6875;
            6876: bcd <= 16'h6876;
            6877: bcd <= 16'h6877;
            6878: bcd <= 16'h6878;
            6879: bcd <= 16'h6879;
            6880: bcd <= 16'h6880;
            6881: bcd <= 16'h6881;
            6882: bcd <= 16'h6882;
            6883: bcd <= 16'h6883;
            6884: bcd <= 16'h6884;
            6885: bcd <= 16'h6885;
            6886: bcd <= 16'h6886;
            6887: bcd <= 16'h6887;
            6888: bcd <= 16'h6888;
            6889: bcd <= 16'h6889;
            6890: bcd <= 16'h6890;
            6891: bcd <= 16'h6891;
            6892: bcd <= 16'h6892;
            6893: bcd <= 16'h6893;
            6894: bcd <= 16'h6894;
            6895: bcd <= 16'h6895;
            6896: bcd <= 16'h6896;
            6897: bcd <= 16'h6897;
            6898: bcd <= 16'h6898;
            6899: bcd <= 16'h6899;
            6900: bcd <= 16'h6900;
            6901: bcd <= 16'h6901;
            6902: bcd <= 16'h6902;
            6903: bcd <= 16'h6903;
            6904: bcd <= 16'h6904;
            6905: bcd <= 16'h6905;
            6906: bcd <= 16'h6906;
            6907: bcd <= 16'h6907;
            6908: bcd <= 16'h6908;
            6909: bcd <= 16'h6909;
            6910: bcd <= 16'h6910;
            6911: bcd <= 16'h6911;
            6912: bcd <= 16'h6912;
            6913: bcd <= 16'h6913;
            6914: bcd <= 16'h6914;
            6915: bcd <= 16'h6915;
            6916: bcd <= 16'h6916;
            6917: bcd <= 16'h6917;
            6918: bcd <= 16'h6918;
            6919: bcd <= 16'h6919;
            6920: bcd <= 16'h6920;
            6921: bcd <= 16'h6921;
            6922: bcd <= 16'h6922;
            6923: bcd <= 16'h6923;
            6924: bcd <= 16'h6924;
            6925: bcd <= 16'h6925;
            6926: bcd <= 16'h6926;
            6927: bcd <= 16'h6927;
            6928: bcd <= 16'h6928;
            6929: bcd <= 16'h6929;
            6930: bcd <= 16'h6930;
            6931: bcd <= 16'h6931;
            6932: bcd <= 16'h6932;
            6933: bcd <= 16'h6933;
            6934: bcd <= 16'h6934;
            6935: bcd <= 16'h6935;
            6936: bcd <= 16'h6936;
            6937: bcd <= 16'h6937;
            6938: bcd <= 16'h6938;
            6939: bcd <= 16'h6939;
            6940: bcd <= 16'h6940;
            6941: bcd <= 16'h6941;
            6942: bcd <= 16'h6942;
            6943: bcd <= 16'h6943;
            6944: bcd <= 16'h6944;
            6945: bcd <= 16'h6945;
            6946: bcd <= 16'h6946;
            6947: bcd <= 16'h6947;
            6948: bcd <= 16'h6948;
            6949: bcd <= 16'h6949;
            6950: bcd <= 16'h6950;
            6951: bcd <= 16'h6951;
            6952: bcd <= 16'h6952;
            6953: bcd <= 16'h6953;
            6954: bcd <= 16'h6954;
            6955: bcd <= 16'h6955;
            6956: bcd <= 16'h6956;
            6957: bcd <= 16'h6957;
            6958: bcd <= 16'h6958;
            6959: bcd <= 16'h6959;
            6960: bcd <= 16'h6960;
            6961: bcd <= 16'h6961;
            6962: bcd <= 16'h6962;
            6963: bcd <= 16'h6963;
            6964: bcd <= 16'h6964;
            6965: bcd <= 16'h6965;
            6966: bcd <= 16'h6966;
            6967: bcd <= 16'h6967;
            6968: bcd <= 16'h6968;
            6969: bcd <= 16'h6969;
            6970: bcd <= 16'h6970;
            6971: bcd <= 16'h6971;
            6972: bcd <= 16'h6972;
            6973: bcd <= 16'h6973;
            6974: bcd <= 16'h6974;
            6975: bcd <= 16'h6975;
            6976: bcd <= 16'h6976;
            6977: bcd <= 16'h6977;
            6978: bcd <= 16'h6978;
            6979: bcd <= 16'h6979;
            6980: bcd <= 16'h6980;
            6981: bcd <= 16'h6981;
            6982: bcd <= 16'h6982;
            6983: bcd <= 16'h6983;
            6984: bcd <= 16'h6984;
            6985: bcd <= 16'h6985;
            6986: bcd <= 16'h6986;
            6987: bcd <= 16'h6987;
            6988: bcd <= 16'h6988;
            6989: bcd <= 16'h6989;
            6990: bcd <= 16'h6990;
            6991: bcd <= 16'h6991;
            6992: bcd <= 16'h6992;
            6993: bcd <= 16'h6993;
            6994: bcd <= 16'h6994;
            6995: bcd <= 16'h6995;
            6996: bcd <= 16'h6996;
            6997: bcd <= 16'h6997;
            6998: bcd <= 16'h6998;
            6999: bcd <= 16'h6999;
            7000: bcd <= 16'h7000;
            7001: bcd <= 16'h7001;
            7002: bcd <= 16'h7002;
            7003: bcd <= 16'h7003;
            7004: bcd <= 16'h7004;
            7005: bcd <= 16'h7005;
            7006: bcd <= 16'h7006;
            7007: bcd <= 16'h7007;
            7008: bcd <= 16'h7008;
            7009: bcd <= 16'h7009;
            7010: bcd <= 16'h7010;
            7011: bcd <= 16'h7011;
            7012: bcd <= 16'h7012;
            7013: bcd <= 16'h7013;
            7014: bcd <= 16'h7014;
            7015: bcd <= 16'h7015;
            7016: bcd <= 16'h7016;
            7017: bcd <= 16'h7017;
            7018: bcd <= 16'h7018;
            7019: bcd <= 16'h7019;
            7020: bcd <= 16'h7020;
            7021: bcd <= 16'h7021;
            7022: bcd <= 16'h7022;
            7023: bcd <= 16'h7023;
            7024: bcd <= 16'h7024;
            7025: bcd <= 16'h7025;
            7026: bcd <= 16'h7026;
            7027: bcd <= 16'h7027;
            7028: bcd <= 16'h7028;
            7029: bcd <= 16'h7029;
            7030: bcd <= 16'h7030;
            7031: bcd <= 16'h7031;
            7032: bcd <= 16'h7032;
            7033: bcd <= 16'h7033;
            7034: bcd <= 16'h7034;
            7035: bcd <= 16'h7035;
            7036: bcd <= 16'h7036;
            7037: bcd <= 16'h7037;
            7038: bcd <= 16'h7038;
            7039: bcd <= 16'h7039;
            7040: bcd <= 16'h7040;
            7041: bcd <= 16'h7041;
            7042: bcd <= 16'h7042;
            7043: bcd <= 16'h7043;
            7044: bcd <= 16'h7044;
            7045: bcd <= 16'h7045;
            7046: bcd <= 16'h7046;
            7047: bcd <= 16'h7047;
            7048: bcd <= 16'h7048;
            7049: bcd <= 16'h7049;
            7050: bcd <= 16'h7050;
            7051: bcd <= 16'h7051;
            7052: bcd <= 16'h7052;
            7053: bcd <= 16'h7053;
            7054: bcd <= 16'h7054;
            7055: bcd <= 16'h7055;
            7056: bcd <= 16'h7056;
            7057: bcd <= 16'h7057;
            7058: bcd <= 16'h7058;
            7059: bcd <= 16'h7059;
            7060: bcd <= 16'h7060;
            7061: bcd <= 16'h7061;
            7062: bcd <= 16'h7062;
            7063: bcd <= 16'h7063;
            7064: bcd <= 16'h7064;
            7065: bcd <= 16'h7065;
            7066: bcd <= 16'h7066;
            7067: bcd <= 16'h7067;
            7068: bcd <= 16'h7068;
            7069: bcd <= 16'h7069;
            7070: bcd <= 16'h7070;
            7071: bcd <= 16'h7071;
            7072: bcd <= 16'h7072;
            7073: bcd <= 16'h7073;
            7074: bcd <= 16'h7074;
            7075: bcd <= 16'h7075;
            7076: bcd <= 16'h7076;
            7077: bcd <= 16'h7077;
            7078: bcd <= 16'h7078;
            7079: bcd <= 16'h7079;
            7080: bcd <= 16'h7080;
            7081: bcd <= 16'h7081;
            7082: bcd <= 16'h7082;
            7083: bcd <= 16'h7083;
            7084: bcd <= 16'h7084;
            7085: bcd <= 16'h7085;
            7086: bcd <= 16'h7086;
            7087: bcd <= 16'h7087;
            7088: bcd <= 16'h7088;
            7089: bcd <= 16'h7089;
            7090: bcd <= 16'h7090;
            7091: bcd <= 16'h7091;
            7092: bcd <= 16'h7092;
            7093: bcd <= 16'h7093;
            7094: bcd <= 16'h7094;
            7095: bcd <= 16'h7095;
            7096: bcd <= 16'h7096;
            7097: bcd <= 16'h7097;
            7098: bcd <= 16'h7098;
            7099: bcd <= 16'h7099;
            7100: bcd <= 16'h7100;
            7101: bcd <= 16'h7101;
            7102: bcd <= 16'h7102;
            7103: bcd <= 16'h7103;
            7104: bcd <= 16'h7104;
            7105: bcd <= 16'h7105;
            7106: bcd <= 16'h7106;
            7107: bcd <= 16'h7107;
            7108: bcd <= 16'h7108;
            7109: bcd <= 16'h7109;
            7110: bcd <= 16'h7110;
            7111: bcd <= 16'h7111;
            7112: bcd <= 16'h7112;
            7113: bcd <= 16'h7113;
            7114: bcd <= 16'h7114;
            7115: bcd <= 16'h7115;
            7116: bcd <= 16'h7116;
            7117: bcd <= 16'h7117;
            7118: bcd <= 16'h7118;
            7119: bcd <= 16'h7119;
            7120: bcd <= 16'h7120;
            7121: bcd <= 16'h7121;
            7122: bcd <= 16'h7122;
            7123: bcd <= 16'h7123;
            7124: bcd <= 16'h7124;
            7125: bcd <= 16'h7125;
            7126: bcd <= 16'h7126;
            7127: bcd <= 16'h7127;
            7128: bcd <= 16'h7128;
            7129: bcd <= 16'h7129;
            7130: bcd <= 16'h7130;
            7131: bcd <= 16'h7131;
            7132: bcd <= 16'h7132;
            7133: bcd <= 16'h7133;
            7134: bcd <= 16'h7134;
            7135: bcd <= 16'h7135;
            7136: bcd <= 16'h7136;
            7137: bcd <= 16'h7137;
            7138: bcd <= 16'h7138;
            7139: bcd <= 16'h7139;
            7140: bcd <= 16'h7140;
            7141: bcd <= 16'h7141;
            7142: bcd <= 16'h7142;
            7143: bcd <= 16'h7143;
            7144: bcd <= 16'h7144;
            7145: bcd <= 16'h7145;
            7146: bcd <= 16'h7146;
            7147: bcd <= 16'h7147;
            7148: bcd <= 16'h7148;
            7149: bcd <= 16'h7149;
            7150: bcd <= 16'h7150;
            7151: bcd <= 16'h7151;
            7152: bcd <= 16'h7152;
            7153: bcd <= 16'h7153;
            7154: bcd <= 16'h7154;
            7155: bcd <= 16'h7155;
            7156: bcd <= 16'h7156;
            7157: bcd <= 16'h7157;
            7158: bcd <= 16'h7158;
            7159: bcd <= 16'h7159;
            7160: bcd <= 16'h7160;
            7161: bcd <= 16'h7161;
            7162: bcd <= 16'h7162;
            7163: bcd <= 16'h7163;
            7164: bcd <= 16'h7164;
            7165: bcd <= 16'h7165;
            7166: bcd <= 16'h7166;
            7167: bcd <= 16'h7167;
            7168: bcd <= 16'h7168;
            7169: bcd <= 16'h7169;
            7170: bcd <= 16'h7170;
            7171: bcd <= 16'h7171;
            7172: bcd <= 16'h7172;
            7173: bcd <= 16'h7173;
            7174: bcd <= 16'h7174;
            7175: bcd <= 16'h7175;
            7176: bcd <= 16'h7176;
            7177: bcd <= 16'h7177;
            7178: bcd <= 16'h7178;
            7179: bcd <= 16'h7179;
            7180: bcd <= 16'h7180;
            7181: bcd <= 16'h7181;
            7182: bcd <= 16'h7182;
            7183: bcd <= 16'h7183;
            7184: bcd <= 16'h7184;
            7185: bcd <= 16'h7185;
            7186: bcd <= 16'h7186;
            7187: bcd <= 16'h7187;
            7188: bcd <= 16'h7188;
            7189: bcd <= 16'h7189;
            7190: bcd <= 16'h7190;
            7191: bcd <= 16'h7191;
            7192: bcd <= 16'h7192;
            7193: bcd <= 16'h7193;
            7194: bcd <= 16'h7194;
            7195: bcd <= 16'h7195;
            7196: bcd <= 16'h7196;
            7197: bcd <= 16'h7197;
            7198: bcd <= 16'h7198;
            7199: bcd <= 16'h7199;
            7200: bcd <= 16'h7200;
            7201: bcd <= 16'h7201;
            7202: bcd <= 16'h7202;
            7203: bcd <= 16'h7203;
            7204: bcd <= 16'h7204;
            7205: bcd <= 16'h7205;
            7206: bcd <= 16'h7206;
            7207: bcd <= 16'h7207;
            7208: bcd <= 16'h7208;
            7209: bcd <= 16'h7209;
            7210: bcd <= 16'h7210;
            7211: bcd <= 16'h7211;
            7212: bcd <= 16'h7212;
            7213: bcd <= 16'h7213;
            7214: bcd <= 16'h7214;
            7215: bcd <= 16'h7215;
            7216: bcd <= 16'h7216;
            7217: bcd <= 16'h7217;
            7218: bcd <= 16'h7218;
            7219: bcd <= 16'h7219;
            7220: bcd <= 16'h7220;
            7221: bcd <= 16'h7221;
            7222: bcd <= 16'h7222;
            7223: bcd <= 16'h7223;
            7224: bcd <= 16'h7224;
            7225: bcd <= 16'h7225;
            7226: bcd <= 16'h7226;
            7227: bcd <= 16'h7227;
            7228: bcd <= 16'h7228;
            7229: bcd <= 16'h7229;
            7230: bcd <= 16'h7230;
            7231: bcd <= 16'h7231;
            7232: bcd <= 16'h7232;
            7233: bcd <= 16'h7233;
            7234: bcd <= 16'h7234;
            7235: bcd <= 16'h7235;
            7236: bcd <= 16'h7236;
            7237: bcd <= 16'h7237;
            7238: bcd <= 16'h7238;
            7239: bcd <= 16'h7239;
            7240: bcd <= 16'h7240;
            7241: bcd <= 16'h7241;
            7242: bcd <= 16'h7242;
            7243: bcd <= 16'h7243;
            7244: bcd <= 16'h7244;
            7245: bcd <= 16'h7245;
            7246: bcd <= 16'h7246;
            7247: bcd <= 16'h7247;
            7248: bcd <= 16'h7248;
            7249: bcd <= 16'h7249;
            7250: bcd <= 16'h7250;
            7251: bcd <= 16'h7251;
            7252: bcd <= 16'h7252;
            7253: bcd <= 16'h7253;
            7254: bcd <= 16'h7254;
            7255: bcd <= 16'h7255;
            7256: bcd <= 16'h7256;
            7257: bcd <= 16'h7257;
            7258: bcd <= 16'h7258;
            7259: bcd <= 16'h7259;
            7260: bcd <= 16'h7260;
            7261: bcd <= 16'h7261;
            7262: bcd <= 16'h7262;
            7263: bcd <= 16'h7263;
            7264: bcd <= 16'h7264;
            7265: bcd <= 16'h7265;
            7266: bcd <= 16'h7266;
            7267: bcd <= 16'h7267;
            7268: bcd <= 16'h7268;
            7269: bcd <= 16'h7269;
            7270: bcd <= 16'h7270;
            7271: bcd <= 16'h7271;
            7272: bcd <= 16'h7272;
            7273: bcd <= 16'h7273;
            7274: bcd <= 16'h7274;
            7275: bcd <= 16'h7275;
            7276: bcd <= 16'h7276;
            7277: bcd <= 16'h7277;
            7278: bcd <= 16'h7278;
            7279: bcd <= 16'h7279;
            7280: bcd <= 16'h7280;
            7281: bcd <= 16'h7281;
            7282: bcd <= 16'h7282;
            7283: bcd <= 16'h7283;
            7284: bcd <= 16'h7284;
            7285: bcd <= 16'h7285;
            7286: bcd <= 16'h7286;
            7287: bcd <= 16'h7287;
            7288: bcd <= 16'h7288;
            7289: bcd <= 16'h7289;
            7290: bcd <= 16'h7290;
            7291: bcd <= 16'h7291;
            7292: bcd <= 16'h7292;
            7293: bcd <= 16'h7293;
            7294: bcd <= 16'h7294;
            7295: bcd <= 16'h7295;
            7296: bcd <= 16'h7296;
            7297: bcd <= 16'h7297;
            7298: bcd <= 16'h7298;
            7299: bcd <= 16'h7299;
            7300: bcd <= 16'h7300;
            7301: bcd <= 16'h7301;
            7302: bcd <= 16'h7302;
            7303: bcd <= 16'h7303;
            7304: bcd <= 16'h7304;
            7305: bcd <= 16'h7305;
            7306: bcd <= 16'h7306;
            7307: bcd <= 16'h7307;
            7308: bcd <= 16'h7308;
            7309: bcd <= 16'h7309;
            7310: bcd <= 16'h7310;
            7311: bcd <= 16'h7311;
            7312: bcd <= 16'h7312;
            7313: bcd <= 16'h7313;
            7314: bcd <= 16'h7314;
            7315: bcd <= 16'h7315;
            7316: bcd <= 16'h7316;
            7317: bcd <= 16'h7317;
            7318: bcd <= 16'h7318;
            7319: bcd <= 16'h7319;
            7320: bcd <= 16'h7320;
            7321: bcd <= 16'h7321;
            7322: bcd <= 16'h7322;
            7323: bcd <= 16'h7323;
            7324: bcd <= 16'h7324;
            7325: bcd <= 16'h7325;
            7326: bcd <= 16'h7326;
            7327: bcd <= 16'h7327;
            7328: bcd <= 16'h7328;
            7329: bcd <= 16'h7329;
            7330: bcd <= 16'h7330;
            7331: bcd <= 16'h7331;
            7332: bcd <= 16'h7332;
            7333: bcd <= 16'h7333;
            7334: bcd <= 16'h7334;
            7335: bcd <= 16'h7335;
            7336: bcd <= 16'h7336;
            7337: bcd <= 16'h7337;
            7338: bcd <= 16'h7338;
            7339: bcd <= 16'h7339;
            7340: bcd <= 16'h7340;
            7341: bcd <= 16'h7341;
            7342: bcd <= 16'h7342;
            7343: bcd <= 16'h7343;
            7344: bcd <= 16'h7344;
            7345: bcd <= 16'h7345;
            7346: bcd <= 16'h7346;
            7347: bcd <= 16'h7347;
            7348: bcd <= 16'h7348;
            7349: bcd <= 16'h7349;
            7350: bcd <= 16'h7350;
            7351: bcd <= 16'h7351;
            7352: bcd <= 16'h7352;
            7353: bcd <= 16'h7353;
            7354: bcd <= 16'h7354;
            7355: bcd <= 16'h7355;
            7356: bcd <= 16'h7356;
            7357: bcd <= 16'h7357;
            7358: bcd <= 16'h7358;
            7359: bcd <= 16'h7359;
            7360: bcd <= 16'h7360;
            7361: bcd <= 16'h7361;
            7362: bcd <= 16'h7362;
            7363: bcd <= 16'h7363;
            7364: bcd <= 16'h7364;
            7365: bcd <= 16'h7365;
            7366: bcd <= 16'h7366;
            7367: bcd <= 16'h7367;
            7368: bcd <= 16'h7368;
            7369: bcd <= 16'h7369;
            7370: bcd <= 16'h7370;
            7371: bcd <= 16'h7371;
            7372: bcd <= 16'h7372;
            7373: bcd <= 16'h7373;
            7374: bcd <= 16'h7374;
            7375: bcd <= 16'h7375;
            7376: bcd <= 16'h7376;
            7377: bcd <= 16'h7377;
            7378: bcd <= 16'h7378;
            7379: bcd <= 16'h7379;
            7380: bcd <= 16'h7380;
            7381: bcd <= 16'h7381;
            7382: bcd <= 16'h7382;
            7383: bcd <= 16'h7383;
            7384: bcd <= 16'h7384;
            7385: bcd <= 16'h7385;
            7386: bcd <= 16'h7386;
            7387: bcd <= 16'h7387;
            7388: bcd <= 16'h7388;
            7389: bcd <= 16'h7389;
            7390: bcd <= 16'h7390;
            7391: bcd <= 16'h7391;
            7392: bcd <= 16'h7392;
            7393: bcd <= 16'h7393;
            7394: bcd <= 16'h7394;
            7395: bcd <= 16'h7395;
            7396: bcd <= 16'h7396;
            7397: bcd <= 16'h7397;
            7398: bcd <= 16'h7398;
            7399: bcd <= 16'h7399;
            7400: bcd <= 16'h7400;
            7401: bcd <= 16'h7401;
            7402: bcd <= 16'h7402;
            7403: bcd <= 16'h7403;
            7404: bcd <= 16'h7404;
            7405: bcd <= 16'h7405;
            7406: bcd <= 16'h7406;
            7407: bcd <= 16'h7407;
            7408: bcd <= 16'h7408;
            7409: bcd <= 16'h7409;
            7410: bcd <= 16'h7410;
            7411: bcd <= 16'h7411;
            7412: bcd <= 16'h7412;
            7413: bcd <= 16'h7413;
            7414: bcd <= 16'h7414;
            7415: bcd <= 16'h7415;
            7416: bcd <= 16'h7416;
            7417: bcd <= 16'h7417;
            7418: bcd <= 16'h7418;
            7419: bcd <= 16'h7419;
            7420: bcd <= 16'h7420;
            7421: bcd <= 16'h7421;
            7422: bcd <= 16'h7422;
            7423: bcd <= 16'h7423;
            7424: bcd <= 16'h7424;
            7425: bcd <= 16'h7425;
            7426: bcd <= 16'h7426;
            7427: bcd <= 16'h7427;
            7428: bcd <= 16'h7428;
            7429: bcd <= 16'h7429;
            7430: bcd <= 16'h7430;
            7431: bcd <= 16'h7431;
            7432: bcd <= 16'h7432;
            7433: bcd <= 16'h7433;
            7434: bcd <= 16'h7434;
            7435: bcd <= 16'h7435;
            7436: bcd <= 16'h7436;
            7437: bcd <= 16'h7437;
            7438: bcd <= 16'h7438;
            7439: bcd <= 16'h7439;
            7440: bcd <= 16'h7440;
            7441: bcd <= 16'h7441;
            7442: bcd <= 16'h7442;
            7443: bcd <= 16'h7443;
            7444: bcd <= 16'h7444;
            7445: bcd <= 16'h7445;
            7446: bcd <= 16'h7446;
            7447: bcd <= 16'h7447;
            7448: bcd <= 16'h7448;
            7449: bcd <= 16'h7449;
            7450: bcd <= 16'h7450;
            7451: bcd <= 16'h7451;
            7452: bcd <= 16'h7452;
            7453: bcd <= 16'h7453;
            7454: bcd <= 16'h7454;
            7455: bcd <= 16'h7455;
            7456: bcd <= 16'h7456;
            7457: bcd <= 16'h7457;
            7458: bcd <= 16'h7458;
            7459: bcd <= 16'h7459;
            7460: bcd <= 16'h7460;
            7461: bcd <= 16'h7461;
            7462: bcd <= 16'h7462;
            7463: bcd <= 16'h7463;
            7464: bcd <= 16'h7464;
            7465: bcd <= 16'h7465;
            7466: bcd <= 16'h7466;
            7467: bcd <= 16'h7467;
            7468: bcd <= 16'h7468;
            7469: bcd <= 16'h7469;
            7470: bcd <= 16'h7470;
            7471: bcd <= 16'h7471;
            7472: bcd <= 16'h7472;
            7473: bcd <= 16'h7473;
            7474: bcd <= 16'h7474;
            7475: bcd <= 16'h7475;
            7476: bcd <= 16'h7476;
            7477: bcd <= 16'h7477;
            7478: bcd <= 16'h7478;
            7479: bcd <= 16'h7479;
            7480: bcd <= 16'h7480;
            7481: bcd <= 16'h7481;
            7482: bcd <= 16'h7482;
            7483: bcd <= 16'h7483;
            7484: bcd <= 16'h7484;
            7485: bcd <= 16'h7485;
            7486: bcd <= 16'h7486;
            7487: bcd <= 16'h7487;
            7488: bcd <= 16'h7488;
            7489: bcd <= 16'h7489;
            7490: bcd <= 16'h7490;
            7491: bcd <= 16'h7491;
            7492: bcd <= 16'h7492;
            7493: bcd <= 16'h7493;
            7494: bcd <= 16'h7494;
            7495: bcd <= 16'h7495;
            7496: bcd <= 16'h7496;
            7497: bcd <= 16'h7497;
            7498: bcd <= 16'h7498;
            7499: bcd <= 16'h7499;
            7500: bcd <= 16'h7500;
            7501: bcd <= 16'h7501;
            7502: bcd <= 16'h7502;
            7503: bcd <= 16'h7503;
            7504: bcd <= 16'h7504;
            7505: bcd <= 16'h7505;
            7506: bcd <= 16'h7506;
            7507: bcd <= 16'h7507;
            7508: bcd <= 16'h7508;
            7509: bcd <= 16'h7509;
            7510: bcd <= 16'h7510;
            7511: bcd <= 16'h7511;
            7512: bcd <= 16'h7512;
            7513: bcd <= 16'h7513;
            7514: bcd <= 16'h7514;
            7515: bcd <= 16'h7515;
            7516: bcd <= 16'h7516;
            7517: bcd <= 16'h7517;
            7518: bcd <= 16'h7518;
            7519: bcd <= 16'h7519;
            7520: bcd <= 16'h7520;
            7521: bcd <= 16'h7521;
            7522: bcd <= 16'h7522;
            7523: bcd <= 16'h7523;
            7524: bcd <= 16'h7524;
            7525: bcd <= 16'h7525;
            7526: bcd <= 16'h7526;
            7527: bcd <= 16'h7527;
            7528: bcd <= 16'h7528;
            7529: bcd <= 16'h7529;
            7530: bcd <= 16'h7530;
            7531: bcd <= 16'h7531;
            7532: bcd <= 16'h7532;
            7533: bcd <= 16'h7533;
            7534: bcd <= 16'h7534;
            7535: bcd <= 16'h7535;
            7536: bcd <= 16'h7536;
            7537: bcd <= 16'h7537;
            7538: bcd <= 16'h7538;
            7539: bcd <= 16'h7539;
            7540: bcd <= 16'h7540;
            7541: bcd <= 16'h7541;
            7542: bcd <= 16'h7542;
            7543: bcd <= 16'h7543;
            7544: bcd <= 16'h7544;
            7545: bcd <= 16'h7545;
            7546: bcd <= 16'h7546;
            7547: bcd <= 16'h7547;
            7548: bcd <= 16'h7548;
            7549: bcd <= 16'h7549;
            7550: bcd <= 16'h7550;
            7551: bcd <= 16'h7551;
            7552: bcd <= 16'h7552;
            7553: bcd <= 16'h7553;
            7554: bcd <= 16'h7554;
            7555: bcd <= 16'h7555;
            7556: bcd <= 16'h7556;
            7557: bcd <= 16'h7557;
            7558: bcd <= 16'h7558;
            7559: bcd <= 16'h7559;
            7560: bcd <= 16'h7560;
            7561: bcd <= 16'h7561;
            7562: bcd <= 16'h7562;
            7563: bcd <= 16'h7563;
            7564: bcd <= 16'h7564;
            7565: bcd <= 16'h7565;
            7566: bcd <= 16'h7566;
            7567: bcd <= 16'h7567;
            7568: bcd <= 16'h7568;
            7569: bcd <= 16'h7569;
            7570: bcd <= 16'h7570;
            7571: bcd <= 16'h7571;
            7572: bcd <= 16'h7572;
            7573: bcd <= 16'h7573;
            7574: bcd <= 16'h7574;
            7575: bcd <= 16'h7575;
            7576: bcd <= 16'h7576;
            7577: bcd <= 16'h7577;
            7578: bcd <= 16'h7578;
            7579: bcd <= 16'h7579;
            7580: bcd <= 16'h7580;
            7581: bcd <= 16'h7581;
            7582: bcd <= 16'h7582;
            7583: bcd <= 16'h7583;
            7584: bcd <= 16'h7584;
            7585: bcd <= 16'h7585;
            7586: bcd <= 16'h7586;
            7587: bcd <= 16'h7587;
            7588: bcd <= 16'h7588;
            7589: bcd <= 16'h7589;
            7590: bcd <= 16'h7590;
            7591: bcd <= 16'h7591;
            7592: bcd <= 16'h7592;
            7593: bcd <= 16'h7593;
            7594: bcd <= 16'h7594;
            7595: bcd <= 16'h7595;
            7596: bcd <= 16'h7596;
            7597: bcd <= 16'h7597;
            7598: bcd <= 16'h7598;
            7599: bcd <= 16'h7599;
            7600: bcd <= 16'h7600;
            7601: bcd <= 16'h7601;
            7602: bcd <= 16'h7602;
            7603: bcd <= 16'h7603;
            7604: bcd <= 16'h7604;
            7605: bcd <= 16'h7605;
            7606: bcd <= 16'h7606;
            7607: bcd <= 16'h7607;
            7608: bcd <= 16'h7608;
            7609: bcd <= 16'h7609;
            7610: bcd <= 16'h7610;
            7611: bcd <= 16'h7611;
            7612: bcd <= 16'h7612;
            7613: bcd <= 16'h7613;
            7614: bcd <= 16'h7614;
            7615: bcd <= 16'h7615;
            7616: bcd <= 16'h7616;
            7617: bcd <= 16'h7617;
            7618: bcd <= 16'h7618;
            7619: bcd <= 16'h7619;
            7620: bcd <= 16'h7620;
            7621: bcd <= 16'h7621;
            7622: bcd <= 16'h7622;
            7623: bcd <= 16'h7623;
            7624: bcd <= 16'h7624;
            7625: bcd <= 16'h7625;
            7626: bcd <= 16'h7626;
            7627: bcd <= 16'h7627;
            7628: bcd <= 16'h7628;
            7629: bcd <= 16'h7629;
            7630: bcd <= 16'h7630;
            7631: bcd <= 16'h7631;
            7632: bcd <= 16'h7632;
            7633: bcd <= 16'h7633;
            7634: bcd <= 16'h7634;
            7635: bcd <= 16'h7635;
            7636: bcd <= 16'h7636;
            7637: bcd <= 16'h7637;
            7638: bcd <= 16'h7638;
            7639: bcd <= 16'h7639;
            7640: bcd <= 16'h7640;
            7641: bcd <= 16'h7641;
            7642: bcd <= 16'h7642;
            7643: bcd <= 16'h7643;
            7644: bcd <= 16'h7644;
            7645: bcd <= 16'h7645;
            7646: bcd <= 16'h7646;
            7647: bcd <= 16'h7647;
            7648: bcd <= 16'h7648;
            7649: bcd <= 16'h7649;
            7650: bcd <= 16'h7650;
            7651: bcd <= 16'h7651;
            7652: bcd <= 16'h7652;
            7653: bcd <= 16'h7653;
            7654: bcd <= 16'h7654;
            7655: bcd <= 16'h7655;
            7656: bcd <= 16'h7656;
            7657: bcd <= 16'h7657;
            7658: bcd <= 16'h7658;
            7659: bcd <= 16'h7659;
            7660: bcd <= 16'h7660;
            7661: bcd <= 16'h7661;
            7662: bcd <= 16'h7662;
            7663: bcd <= 16'h7663;
            7664: bcd <= 16'h7664;
            7665: bcd <= 16'h7665;
            7666: bcd <= 16'h7666;
            7667: bcd <= 16'h7667;
            7668: bcd <= 16'h7668;
            7669: bcd <= 16'h7669;
            7670: bcd <= 16'h7670;
            7671: bcd <= 16'h7671;
            7672: bcd <= 16'h7672;
            7673: bcd <= 16'h7673;
            7674: bcd <= 16'h7674;
            7675: bcd <= 16'h7675;
            7676: bcd <= 16'h7676;
            7677: bcd <= 16'h7677;
            7678: bcd <= 16'h7678;
            7679: bcd <= 16'h7679;
            7680: bcd <= 16'h7680;
            7681: bcd <= 16'h7681;
            7682: bcd <= 16'h7682;
            7683: bcd <= 16'h7683;
            7684: bcd <= 16'h7684;
            7685: bcd <= 16'h7685;
            7686: bcd <= 16'h7686;
            7687: bcd <= 16'h7687;
            7688: bcd <= 16'h7688;
            7689: bcd <= 16'h7689;
            7690: bcd <= 16'h7690;
            7691: bcd <= 16'h7691;
            7692: bcd <= 16'h7692;
            7693: bcd <= 16'h7693;
            7694: bcd <= 16'h7694;
            7695: bcd <= 16'h7695;
            7696: bcd <= 16'h7696;
            7697: bcd <= 16'h7697;
            7698: bcd <= 16'h7698;
            7699: bcd <= 16'h7699;
            7700: bcd <= 16'h7700;
            7701: bcd <= 16'h7701;
            7702: bcd <= 16'h7702;
            7703: bcd <= 16'h7703;
            7704: bcd <= 16'h7704;
            7705: bcd <= 16'h7705;
            7706: bcd <= 16'h7706;
            7707: bcd <= 16'h7707;
            7708: bcd <= 16'h7708;
            7709: bcd <= 16'h7709;
            7710: bcd <= 16'h7710;
            7711: bcd <= 16'h7711;
            7712: bcd <= 16'h7712;
            7713: bcd <= 16'h7713;
            7714: bcd <= 16'h7714;
            7715: bcd <= 16'h7715;
            7716: bcd <= 16'h7716;
            7717: bcd <= 16'h7717;
            7718: bcd <= 16'h7718;
            7719: bcd <= 16'h7719;
            7720: bcd <= 16'h7720;
            7721: bcd <= 16'h7721;
            7722: bcd <= 16'h7722;
            7723: bcd <= 16'h7723;
            7724: bcd <= 16'h7724;
            7725: bcd <= 16'h7725;
            7726: bcd <= 16'h7726;
            7727: bcd <= 16'h7727;
            7728: bcd <= 16'h7728;
            7729: bcd <= 16'h7729;
            7730: bcd <= 16'h7730;
            7731: bcd <= 16'h7731;
            7732: bcd <= 16'h7732;
            7733: bcd <= 16'h7733;
            7734: bcd <= 16'h7734;
            7735: bcd <= 16'h7735;
            7736: bcd <= 16'h7736;
            7737: bcd <= 16'h7737;
            7738: bcd <= 16'h7738;
            7739: bcd <= 16'h7739;
            7740: bcd <= 16'h7740;
            7741: bcd <= 16'h7741;
            7742: bcd <= 16'h7742;
            7743: bcd <= 16'h7743;
            7744: bcd <= 16'h7744;
            7745: bcd <= 16'h7745;
            7746: bcd <= 16'h7746;
            7747: bcd <= 16'h7747;
            7748: bcd <= 16'h7748;
            7749: bcd <= 16'h7749;
            7750: bcd <= 16'h7750;
            7751: bcd <= 16'h7751;
            7752: bcd <= 16'h7752;
            7753: bcd <= 16'h7753;
            7754: bcd <= 16'h7754;
            7755: bcd <= 16'h7755;
            7756: bcd <= 16'h7756;
            7757: bcd <= 16'h7757;
            7758: bcd <= 16'h7758;
            7759: bcd <= 16'h7759;
            7760: bcd <= 16'h7760;
            7761: bcd <= 16'h7761;
            7762: bcd <= 16'h7762;
            7763: bcd <= 16'h7763;
            7764: bcd <= 16'h7764;
            7765: bcd <= 16'h7765;
            7766: bcd <= 16'h7766;
            7767: bcd <= 16'h7767;
            7768: bcd <= 16'h7768;
            7769: bcd <= 16'h7769;
            7770: bcd <= 16'h7770;
            7771: bcd <= 16'h7771;
            7772: bcd <= 16'h7772;
            7773: bcd <= 16'h7773;
            7774: bcd <= 16'h7774;
            7775: bcd <= 16'h7775;
            7776: bcd <= 16'h7776;
            7777: bcd <= 16'h7777;
            7778: bcd <= 16'h7778;
            7779: bcd <= 16'h7779;
            7780: bcd <= 16'h7780;
            7781: bcd <= 16'h7781;
            7782: bcd <= 16'h7782;
            7783: bcd <= 16'h7783;
            7784: bcd <= 16'h7784;
            7785: bcd <= 16'h7785;
            7786: bcd <= 16'h7786;
            7787: bcd <= 16'h7787;
            7788: bcd <= 16'h7788;
            7789: bcd <= 16'h7789;
            7790: bcd <= 16'h7790;
            7791: bcd <= 16'h7791;
            7792: bcd <= 16'h7792;
            7793: bcd <= 16'h7793;
            7794: bcd <= 16'h7794;
            7795: bcd <= 16'h7795;
            7796: bcd <= 16'h7796;
            7797: bcd <= 16'h7797;
            7798: bcd <= 16'h7798;
            7799: bcd <= 16'h7799;
            7800: bcd <= 16'h7800;
            7801: bcd <= 16'h7801;
            7802: bcd <= 16'h7802;
            7803: bcd <= 16'h7803;
            7804: bcd <= 16'h7804;
            7805: bcd <= 16'h7805;
            7806: bcd <= 16'h7806;
            7807: bcd <= 16'h7807;
            7808: bcd <= 16'h7808;
            7809: bcd <= 16'h7809;
            7810: bcd <= 16'h7810;
            7811: bcd <= 16'h7811;
            7812: bcd <= 16'h7812;
            7813: bcd <= 16'h7813;
            7814: bcd <= 16'h7814;
            7815: bcd <= 16'h7815;
            7816: bcd <= 16'h7816;
            7817: bcd <= 16'h7817;
            7818: bcd <= 16'h7818;
            7819: bcd <= 16'h7819;
            7820: bcd <= 16'h7820;
            7821: bcd <= 16'h7821;
            7822: bcd <= 16'h7822;
            7823: bcd <= 16'h7823;
            7824: bcd <= 16'h7824;
            7825: bcd <= 16'h7825;
            7826: bcd <= 16'h7826;
            7827: bcd <= 16'h7827;
            7828: bcd <= 16'h7828;
            7829: bcd <= 16'h7829;
            7830: bcd <= 16'h7830;
            7831: bcd <= 16'h7831;
            7832: bcd <= 16'h7832;
            7833: bcd <= 16'h7833;
            7834: bcd <= 16'h7834;
            7835: bcd <= 16'h7835;
            7836: bcd <= 16'h7836;
            7837: bcd <= 16'h7837;
            7838: bcd <= 16'h7838;
            7839: bcd <= 16'h7839;
            7840: bcd <= 16'h7840;
            7841: bcd <= 16'h7841;
            7842: bcd <= 16'h7842;
            7843: bcd <= 16'h7843;
            7844: bcd <= 16'h7844;
            7845: bcd <= 16'h7845;
            7846: bcd <= 16'h7846;
            7847: bcd <= 16'h7847;
            7848: bcd <= 16'h7848;
            7849: bcd <= 16'h7849;
            7850: bcd <= 16'h7850;
            7851: bcd <= 16'h7851;
            7852: bcd <= 16'h7852;
            7853: bcd <= 16'h7853;
            7854: bcd <= 16'h7854;
            7855: bcd <= 16'h7855;
            7856: bcd <= 16'h7856;
            7857: bcd <= 16'h7857;
            7858: bcd <= 16'h7858;
            7859: bcd <= 16'h7859;
            7860: bcd <= 16'h7860;
            7861: bcd <= 16'h7861;
            7862: bcd <= 16'h7862;
            7863: bcd <= 16'h7863;
            7864: bcd <= 16'h7864;
            7865: bcd <= 16'h7865;
            7866: bcd <= 16'h7866;
            7867: bcd <= 16'h7867;
            7868: bcd <= 16'h7868;
            7869: bcd <= 16'h7869;
            7870: bcd <= 16'h7870;
            7871: bcd <= 16'h7871;
            7872: bcd <= 16'h7872;
            7873: bcd <= 16'h7873;
            7874: bcd <= 16'h7874;
            7875: bcd <= 16'h7875;
            7876: bcd <= 16'h7876;
            7877: bcd <= 16'h7877;
            7878: bcd <= 16'h7878;
            7879: bcd <= 16'h7879;
            7880: bcd <= 16'h7880;
            7881: bcd <= 16'h7881;
            7882: bcd <= 16'h7882;
            7883: bcd <= 16'h7883;
            7884: bcd <= 16'h7884;
            7885: bcd <= 16'h7885;
            7886: bcd <= 16'h7886;
            7887: bcd <= 16'h7887;
            7888: bcd <= 16'h7888;
            7889: bcd <= 16'h7889;
            7890: bcd <= 16'h7890;
            7891: bcd <= 16'h7891;
            7892: bcd <= 16'h7892;
            7893: bcd <= 16'h7893;
            7894: bcd <= 16'h7894;
            7895: bcd <= 16'h7895;
            7896: bcd <= 16'h7896;
            7897: bcd <= 16'h7897;
            7898: bcd <= 16'h7898;
            7899: bcd <= 16'h7899;
            7900: bcd <= 16'h7900;
            7901: bcd <= 16'h7901;
            7902: bcd <= 16'h7902;
            7903: bcd <= 16'h7903;
            7904: bcd <= 16'h7904;
            7905: bcd <= 16'h7905;
            7906: bcd <= 16'h7906;
            7907: bcd <= 16'h7907;
            7908: bcd <= 16'h7908;
            7909: bcd <= 16'h7909;
            7910: bcd <= 16'h7910;
            7911: bcd <= 16'h7911;
            7912: bcd <= 16'h7912;
            7913: bcd <= 16'h7913;
            7914: bcd <= 16'h7914;
            7915: bcd <= 16'h7915;
            7916: bcd <= 16'h7916;
            7917: bcd <= 16'h7917;
            7918: bcd <= 16'h7918;
            7919: bcd <= 16'h7919;
            7920: bcd <= 16'h7920;
            7921: bcd <= 16'h7921;
            7922: bcd <= 16'h7922;
            7923: bcd <= 16'h7923;
            7924: bcd <= 16'h7924;
            7925: bcd <= 16'h7925;
            7926: bcd <= 16'h7926;
            7927: bcd <= 16'h7927;
            7928: bcd <= 16'h7928;
            7929: bcd <= 16'h7929;
            7930: bcd <= 16'h7930;
            7931: bcd <= 16'h7931;
            7932: bcd <= 16'h7932;
            7933: bcd <= 16'h7933;
            7934: bcd <= 16'h7934;
            7935: bcd <= 16'h7935;
            7936: bcd <= 16'h7936;
            7937: bcd <= 16'h7937;
            7938: bcd <= 16'h7938;
            7939: bcd <= 16'h7939;
            7940: bcd <= 16'h7940;
            7941: bcd <= 16'h7941;
            7942: bcd <= 16'h7942;
            7943: bcd <= 16'h7943;
            7944: bcd <= 16'h7944;
            7945: bcd <= 16'h7945;
            7946: bcd <= 16'h7946;
            7947: bcd <= 16'h7947;
            7948: bcd <= 16'h7948;
            7949: bcd <= 16'h7949;
            7950: bcd <= 16'h7950;
            7951: bcd <= 16'h7951;
            7952: bcd <= 16'h7952;
            7953: bcd <= 16'h7953;
            7954: bcd <= 16'h7954;
            7955: bcd <= 16'h7955;
            7956: bcd <= 16'h7956;
            7957: bcd <= 16'h7957;
            7958: bcd <= 16'h7958;
            7959: bcd <= 16'h7959;
            7960: bcd <= 16'h7960;
            7961: bcd <= 16'h7961;
            7962: bcd <= 16'h7962;
            7963: bcd <= 16'h7963;
            7964: bcd <= 16'h7964;
            7965: bcd <= 16'h7965;
            7966: bcd <= 16'h7966;
            7967: bcd <= 16'h7967;
            7968: bcd <= 16'h7968;
            7969: bcd <= 16'h7969;
            7970: bcd <= 16'h7970;
            7971: bcd <= 16'h7971;
            7972: bcd <= 16'h7972;
            7973: bcd <= 16'h7973;
            7974: bcd <= 16'h7974;
            7975: bcd <= 16'h7975;
            7976: bcd <= 16'h7976;
            7977: bcd <= 16'h7977;
            7978: bcd <= 16'h7978;
            7979: bcd <= 16'h7979;
            7980: bcd <= 16'h7980;
            7981: bcd <= 16'h7981;
            7982: bcd <= 16'h7982;
            7983: bcd <= 16'h7983;
            7984: bcd <= 16'h7984;
            7985: bcd <= 16'h7985;
            7986: bcd <= 16'h7986;
            7987: bcd <= 16'h7987;
            7988: bcd <= 16'h7988;
            7989: bcd <= 16'h7989;
            7990: bcd <= 16'h7990;
            7991: bcd <= 16'h7991;
            7992: bcd <= 16'h7992;
            7993: bcd <= 16'h7993;
            7994: bcd <= 16'h7994;
            7995: bcd <= 16'h7995;
            7996: bcd <= 16'h7996;
            7997: bcd <= 16'h7997;
            7998: bcd <= 16'h7998;
            7999: bcd <= 16'h7999;
            8000: bcd <= 16'h8000;
            8001: bcd <= 16'h8001;
            8002: bcd <= 16'h8002;
            8003: bcd <= 16'h8003;
            8004: bcd <= 16'h8004;
            8005: bcd <= 16'h8005;
            8006: bcd <= 16'h8006;
            8007: bcd <= 16'h8007;
            8008: bcd <= 16'h8008;
            8009: bcd <= 16'h8009;
            8010: bcd <= 16'h8010;
            8011: bcd <= 16'h8011;
            8012: bcd <= 16'h8012;
            8013: bcd <= 16'h8013;
            8014: bcd <= 16'h8014;
            8015: bcd <= 16'h8015;
            8016: bcd <= 16'h8016;
            8017: bcd <= 16'h8017;
            8018: bcd <= 16'h8018;
            8019: bcd <= 16'h8019;
            8020: bcd <= 16'h8020;
            8021: bcd <= 16'h8021;
            8022: bcd <= 16'h8022;
            8023: bcd <= 16'h8023;
            8024: bcd <= 16'h8024;
            8025: bcd <= 16'h8025;
            8026: bcd <= 16'h8026;
            8027: bcd <= 16'h8027;
            8028: bcd <= 16'h8028;
            8029: bcd <= 16'h8029;
            8030: bcd <= 16'h8030;
            8031: bcd <= 16'h8031;
            8032: bcd <= 16'h8032;
            8033: bcd <= 16'h8033;
            8034: bcd <= 16'h8034;
            8035: bcd <= 16'h8035;
            8036: bcd <= 16'h8036;
            8037: bcd <= 16'h8037;
            8038: bcd <= 16'h8038;
            8039: bcd <= 16'h8039;
            8040: bcd <= 16'h8040;
            8041: bcd <= 16'h8041;
            8042: bcd <= 16'h8042;
            8043: bcd <= 16'h8043;
            8044: bcd <= 16'h8044;
            8045: bcd <= 16'h8045;
            8046: bcd <= 16'h8046;
            8047: bcd <= 16'h8047;
            8048: bcd <= 16'h8048;
            8049: bcd <= 16'h8049;
            8050: bcd <= 16'h8050;
            8051: bcd <= 16'h8051;
            8052: bcd <= 16'h8052;
            8053: bcd <= 16'h8053;
            8054: bcd <= 16'h8054;
            8055: bcd <= 16'h8055;
            8056: bcd <= 16'h8056;
            8057: bcd <= 16'h8057;
            8058: bcd <= 16'h8058;
            8059: bcd <= 16'h8059;
            8060: bcd <= 16'h8060;
            8061: bcd <= 16'h8061;
            8062: bcd <= 16'h8062;
            8063: bcd <= 16'h8063;
            8064: bcd <= 16'h8064;
            8065: bcd <= 16'h8065;
            8066: bcd <= 16'h8066;
            8067: bcd <= 16'h8067;
            8068: bcd <= 16'h8068;
            8069: bcd <= 16'h8069;
            8070: bcd <= 16'h8070;
            8071: bcd <= 16'h8071;
            8072: bcd <= 16'h8072;
            8073: bcd <= 16'h8073;
            8074: bcd <= 16'h8074;
            8075: bcd <= 16'h8075;
            8076: bcd <= 16'h8076;
            8077: bcd <= 16'h8077;
            8078: bcd <= 16'h8078;
            8079: bcd <= 16'h8079;
            8080: bcd <= 16'h8080;
            8081: bcd <= 16'h8081;
            8082: bcd <= 16'h8082;
            8083: bcd <= 16'h8083;
            8084: bcd <= 16'h8084;
            8085: bcd <= 16'h8085;
            8086: bcd <= 16'h8086;
            8087: bcd <= 16'h8087;
            8088: bcd <= 16'h8088;
            8089: bcd <= 16'h8089;
            8090: bcd <= 16'h8090;
            8091: bcd <= 16'h8091;
            8092: bcd <= 16'h8092;
            8093: bcd <= 16'h8093;
            8094: bcd <= 16'h8094;
            8095: bcd <= 16'h8095;
            8096: bcd <= 16'h8096;
            8097: bcd <= 16'h8097;
            8098: bcd <= 16'h8098;
            8099: bcd <= 16'h8099;
            8100: bcd <= 16'h8100;
            8101: bcd <= 16'h8101;
            8102: bcd <= 16'h8102;
            8103: bcd <= 16'h8103;
            8104: bcd <= 16'h8104;
            8105: bcd <= 16'h8105;
            8106: bcd <= 16'h8106;
            8107: bcd <= 16'h8107;
            8108: bcd <= 16'h8108;
            8109: bcd <= 16'h8109;
            8110: bcd <= 16'h8110;
            8111: bcd <= 16'h8111;
            8112: bcd <= 16'h8112;
            8113: bcd <= 16'h8113;
            8114: bcd <= 16'h8114;
            8115: bcd <= 16'h8115;
            8116: bcd <= 16'h8116;
            8117: bcd <= 16'h8117;
            8118: bcd <= 16'h8118;
            8119: bcd <= 16'h8119;
            8120: bcd <= 16'h8120;
            8121: bcd <= 16'h8121;
            8122: bcd <= 16'h8122;
            8123: bcd <= 16'h8123;
            8124: bcd <= 16'h8124;
            8125: bcd <= 16'h8125;
            8126: bcd <= 16'h8126;
            8127: bcd <= 16'h8127;
            8128: bcd <= 16'h8128;
            8129: bcd <= 16'h8129;
            8130: bcd <= 16'h8130;
            8131: bcd <= 16'h8131;
            8132: bcd <= 16'h8132;
            8133: bcd <= 16'h8133;
            8134: bcd <= 16'h8134;
            8135: bcd <= 16'h8135;
            8136: bcd <= 16'h8136;
            8137: bcd <= 16'h8137;
            8138: bcd <= 16'h8138;
            8139: bcd <= 16'h8139;
            8140: bcd <= 16'h8140;
            8141: bcd <= 16'h8141;
            8142: bcd <= 16'h8142;
            8143: bcd <= 16'h8143;
            8144: bcd <= 16'h8144;
            8145: bcd <= 16'h8145;
            8146: bcd <= 16'h8146;
            8147: bcd <= 16'h8147;
            8148: bcd <= 16'h8148;
            8149: bcd <= 16'h8149;
            8150: bcd <= 16'h8150;
            8151: bcd <= 16'h8151;
            8152: bcd <= 16'h8152;
            8153: bcd <= 16'h8153;
            8154: bcd <= 16'h8154;
            8155: bcd <= 16'h8155;
            8156: bcd <= 16'h8156;
            8157: bcd <= 16'h8157;
            8158: bcd <= 16'h8158;
            8159: bcd <= 16'h8159;
            8160: bcd <= 16'h8160;
            8161: bcd <= 16'h8161;
            8162: bcd <= 16'h8162;
            8163: bcd <= 16'h8163;
            8164: bcd <= 16'h8164;
            8165: bcd <= 16'h8165;
            8166: bcd <= 16'h8166;
            8167: bcd <= 16'h8167;
            8168: bcd <= 16'h8168;
            8169: bcd <= 16'h8169;
            8170: bcd <= 16'h8170;
            8171: bcd <= 16'h8171;
            8172: bcd <= 16'h8172;
            8173: bcd <= 16'h8173;
            8174: bcd <= 16'h8174;
            8175: bcd <= 16'h8175;
            8176: bcd <= 16'h8176;
            8177: bcd <= 16'h8177;
            8178: bcd <= 16'h8178;
            8179: bcd <= 16'h8179;
            8180: bcd <= 16'h8180;
            8181: bcd <= 16'h8181;
            8182: bcd <= 16'h8182;
            8183: bcd <= 16'h8183;
            8184: bcd <= 16'h8184;
            8185: bcd <= 16'h8185;
            8186: bcd <= 16'h8186;
            8187: bcd <= 16'h8187;
            8188: bcd <= 16'h8188;
            8189: bcd <= 16'h8189;
            8190: bcd <= 16'h8190;
            8191: bcd <= 16'h8191;
            8192: bcd <= 16'h8192;
            8193: bcd <= 16'h8193;
            8194: bcd <= 16'h8194;
            8195: bcd <= 16'h8195;
            8196: bcd <= 16'h8196;
            8197: bcd <= 16'h8197;
            8198: bcd <= 16'h8198;
            8199: bcd <= 16'h8199;
            8200: bcd <= 16'h8200;
            8201: bcd <= 16'h8201;
            8202: bcd <= 16'h8202;
            8203: bcd <= 16'h8203;
            8204: bcd <= 16'h8204;
            8205: bcd <= 16'h8205;
            8206: bcd <= 16'h8206;
            8207: bcd <= 16'h8207;
            8208: bcd <= 16'h8208;
            8209: bcd <= 16'h8209;
            8210: bcd <= 16'h8210;
            8211: bcd <= 16'h8211;
            8212: bcd <= 16'h8212;
            8213: bcd <= 16'h8213;
            8214: bcd <= 16'h8214;
            8215: bcd <= 16'h8215;
            8216: bcd <= 16'h8216;
            8217: bcd <= 16'h8217;
            8218: bcd <= 16'h8218;
            8219: bcd <= 16'h8219;
            8220: bcd <= 16'h8220;
            8221: bcd <= 16'h8221;
            8222: bcd <= 16'h8222;
            8223: bcd <= 16'h8223;
            8224: bcd <= 16'h8224;
            8225: bcd <= 16'h8225;
            8226: bcd <= 16'h8226;
            8227: bcd <= 16'h8227;
            8228: bcd <= 16'h8228;
            8229: bcd <= 16'h8229;
            8230: bcd <= 16'h8230;
            8231: bcd <= 16'h8231;
            8232: bcd <= 16'h8232;
            8233: bcd <= 16'h8233;
            8234: bcd <= 16'h8234;
            8235: bcd <= 16'h8235;
            8236: bcd <= 16'h8236;
            8237: bcd <= 16'h8237;
            8238: bcd <= 16'h8238;
            8239: bcd <= 16'h8239;
            8240: bcd <= 16'h8240;
            8241: bcd <= 16'h8241;
            8242: bcd <= 16'h8242;
            8243: bcd <= 16'h8243;
            8244: bcd <= 16'h8244;
            8245: bcd <= 16'h8245;
            8246: bcd <= 16'h8246;
            8247: bcd <= 16'h8247;
            8248: bcd <= 16'h8248;
            8249: bcd <= 16'h8249;
            8250: bcd <= 16'h8250;
            8251: bcd <= 16'h8251;
            8252: bcd <= 16'h8252;
            8253: bcd <= 16'h8253;
            8254: bcd <= 16'h8254;
            8255: bcd <= 16'h8255;
            8256: bcd <= 16'h8256;
            8257: bcd <= 16'h8257;
            8258: bcd <= 16'h8258;
            8259: bcd <= 16'h8259;
            8260: bcd <= 16'h8260;
            8261: bcd <= 16'h8261;
            8262: bcd <= 16'h8262;
            8263: bcd <= 16'h8263;
            8264: bcd <= 16'h8264;
            8265: bcd <= 16'h8265;
            8266: bcd <= 16'h8266;
            8267: bcd <= 16'h8267;
            8268: bcd <= 16'h8268;
            8269: bcd <= 16'h8269;
            8270: bcd <= 16'h8270;
            8271: bcd <= 16'h8271;
            8272: bcd <= 16'h8272;
            8273: bcd <= 16'h8273;
            8274: bcd <= 16'h8274;
            8275: bcd <= 16'h8275;
            8276: bcd <= 16'h8276;
            8277: bcd <= 16'h8277;
            8278: bcd <= 16'h8278;
            8279: bcd <= 16'h8279;
            8280: bcd <= 16'h8280;
            8281: bcd <= 16'h8281;
            8282: bcd <= 16'h8282;
            8283: bcd <= 16'h8283;
            8284: bcd <= 16'h8284;
            8285: bcd <= 16'h8285;
            8286: bcd <= 16'h8286;
            8287: bcd <= 16'h8287;
            8288: bcd <= 16'h8288;
            8289: bcd <= 16'h8289;
            8290: bcd <= 16'h8290;
            8291: bcd <= 16'h8291;
            8292: bcd <= 16'h8292;
            8293: bcd <= 16'h8293;
            8294: bcd <= 16'h8294;
            8295: bcd <= 16'h8295;
            8296: bcd <= 16'h8296;
            8297: bcd <= 16'h8297;
            8298: bcd <= 16'h8298;
            8299: bcd <= 16'h8299;
            8300: bcd <= 16'h8300;
            8301: bcd <= 16'h8301;
            8302: bcd <= 16'h8302;
            8303: bcd <= 16'h8303;
            8304: bcd <= 16'h8304;
            8305: bcd <= 16'h8305;
            8306: bcd <= 16'h8306;
            8307: bcd <= 16'h8307;
            8308: bcd <= 16'h8308;
            8309: bcd <= 16'h8309;
            8310: bcd <= 16'h8310;
            8311: bcd <= 16'h8311;
            8312: bcd <= 16'h8312;
            8313: bcd <= 16'h8313;
            8314: bcd <= 16'h8314;
            8315: bcd <= 16'h8315;
            8316: bcd <= 16'h8316;
            8317: bcd <= 16'h8317;
            8318: bcd <= 16'h8318;
            8319: bcd <= 16'h8319;
            8320: bcd <= 16'h8320;
            8321: bcd <= 16'h8321;
            8322: bcd <= 16'h8322;
            8323: bcd <= 16'h8323;
            8324: bcd <= 16'h8324;
            8325: bcd <= 16'h8325;
            8326: bcd <= 16'h8326;
            8327: bcd <= 16'h8327;
            8328: bcd <= 16'h8328;
            8329: bcd <= 16'h8329;
            8330: bcd <= 16'h8330;
            8331: bcd <= 16'h8331;
            8332: bcd <= 16'h8332;
            8333: bcd <= 16'h8333;
            8334: bcd <= 16'h8334;
            8335: bcd <= 16'h8335;
            8336: bcd <= 16'h8336;
            8337: bcd <= 16'h8337;
            8338: bcd <= 16'h8338;
            8339: bcd <= 16'h8339;
            8340: bcd <= 16'h8340;
            8341: bcd <= 16'h8341;
            8342: bcd <= 16'h8342;
            8343: bcd <= 16'h8343;
            8344: bcd <= 16'h8344;
            8345: bcd <= 16'h8345;
            8346: bcd <= 16'h8346;
            8347: bcd <= 16'h8347;
            8348: bcd <= 16'h8348;
            8349: bcd <= 16'h8349;
            8350: bcd <= 16'h8350;
            8351: bcd <= 16'h8351;
            8352: bcd <= 16'h8352;
            8353: bcd <= 16'h8353;
            8354: bcd <= 16'h8354;
            8355: bcd <= 16'h8355;
            8356: bcd <= 16'h8356;
            8357: bcd <= 16'h8357;
            8358: bcd <= 16'h8358;
            8359: bcd <= 16'h8359;
            8360: bcd <= 16'h8360;
            8361: bcd <= 16'h8361;
            8362: bcd <= 16'h8362;
            8363: bcd <= 16'h8363;
            8364: bcd <= 16'h8364;
            8365: bcd <= 16'h8365;
            8366: bcd <= 16'h8366;
            8367: bcd <= 16'h8367;
            8368: bcd <= 16'h8368;
            8369: bcd <= 16'h8369;
            8370: bcd <= 16'h8370;
            8371: bcd <= 16'h8371;
            8372: bcd <= 16'h8372;
            8373: bcd <= 16'h8373;
            8374: bcd <= 16'h8374;
            8375: bcd <= 16'h8375;
            8376: bcd <= 16'h8376;
            8377: bcd <= 16'h8377;
            8378: bcd <= 16'h8378;
            8379: bcd <= 16'h8379;
            8380: bcd <= 16'h8380;
            8381: bcd <= 16'h8381;
            8382: bcd <= 16'h8382;
            8383: bcd <= 16'h8383;
            8384: bcd <= 16'h8384;
            8385: bcd <= 16'h8385;
            8386: bcd <= 16'h8386;
            8387: bcd <= 16'h8387;
            8388: bcd <= 16'h8388;
            8389: bcd <= 16'h8389;
            8390: bcd <= 16'h8390;
            8391: bcd <= 16'h8391;
            8392: bcd <= 16'h8392;
            8393: bcd <= 16'h8393;
            8394: bcd <= 16'h8394;
            8395: bcd <= 16'h8395;
            8396: bcd <= 16'h8396;
            8397: bcd <= 16'h8397;
            8398: bcd <= 16'h8398;
            8399: bcd <= 16'h8399;
            8400: bcd <= 16'h8400;
            8401: bcd <= 16'h8401;
            8402: bcd <= 16'h8402;
            8403: bcd <= 16'h8403;
            8404: bcd <= 16'h8404;
            8405: bcd <= 16'h8405;
            8406: bcd <= 16'h8406;
            8407: bcd <= 16'h8407;
            8408: bcd <= 16'h8408;
            8409: bcd <= 16'h8409;
            8410: bcd <= 16'h8410;
            8411: bcd <= 16'h8411;
            8412: bcd <= 16'h8412;
            8413: bcd <= 16'h8413;
            8414: bcd <= 16'h8414;
            8415: bcd <= 16'h8415;
            8416: bcd <= 16'h8416;
            8417: bcd <= 16'h8417;
            8418: bcd <= 16'h8418;
            8419: bcd <= 16'h8419;
            8420: bcd <= 16'h8420;
            8421: bcd <= 16'h8421;
            8422: bcd <= 16'h8422;
            8423: bcd <= 16'h8423;
            8424: bcd <= 16'h8424;
            8425: bcd <= 16'h8425;
            8426: bcd <= 16'h8426;
            8427: bcd <= 16'h8427;
            8428: bcd <= 16'h8428;
            8429: bcd <= 16'h8429;
            8430: bcd <= 16'h8430;
            8431: bcd <= 16'h8431;
            8432: bcd <= 16'h8432;
            8433: bcd <= 16'h8433;
            8434: bcd <= 16'h8434;
            8435: bcd <= 16'h8435;
            8436: bcd <= 16'h8436;
            8437: bcd <= 16'h8437;
            8438: bcd <= 16'h8438;
            8439: bcd <= 16'h8439;
            8440: bcd <= 16'h8440;
            8441: bcd <= 16'h8441;
            8442: bcd <= 16'h8442;
            8443: bcd <= 16'h8443;
            8444: bcd <= 16'h8444;
            8445: bcd <= 16'h8445;
            8446: bcd <= 16'h8446;
            8447: bcd <= 16'h8447;
            8448: bcd <= 16'h8448;
            8449: bcd <= 16'h8449;
            8450: bcd <= 16'h8450;
            8451: bcd <= 16'h8451;
            8452: bcd <= 16'h8452;
            8453: bcd <= 16'h8453;
            8454: bcd <= 16'h8454;
            8455: bcd <= 16'h8455;
            8456: bcd <= 16'h8456;
            8457: bcd <= 16'h8457;
            8458: bcd <= 16'h8458;
            8459: bcd <= 16'h8459;
            8460: bcd <= 16'h8460;
            8461: bcd <= 16'h8461;
            8462: bcd <= 16'h8462;
            8463: bcd <= 16'h8463;
            8464: bcd <= 16'h8464;
            8465: bcd <= 16'h8465;
            8466: bcd <= 16'h8466;
            8467: bcd <= 16'h8467;
            8468: bcd <= 16'h8468;
            8469: bcd <= 16'h8469;
            8470: bcd <= 16'h8470;
            8471: bcd <= 16'h8471;
            8472: bcd <= 16'h8472;
            8473: bcd <= 16'h8473;
            8474: bcd <= 16'h8474;
            8475: bcd <= 16'h8475;
            8476: bcd <= 16'h8476;
            8477: bcd <= 16'h8477;
            8478: bcd <= 16'h8478;
            8479: bcd <= 16'h8479;
            8480: bcd <= 16'h8480;
            8481: bcd <= 16'h8481;
            8482: bcd <= 16'h8482;
            8483: bcd <= 16'h8483;
            8484: bcd <= 16'h8484;
            8485: bcd <= 16'h8485;
            8486: bcd <= 16'h8486;
            8487: bcd <= 16'h8487;
            8488: bcd <= 16'h8488;
            8489: bcd <= 16'h8489;
            8490: bcd <= 16'h8490;
            8491: bcd <= 16'h8491;
            8492: bcd <= 16'h8492;
            8493: bcd <= 16'h8493;
            8494: bcd <= 16'h8494;
            8495: bcd <= 16'h8495;
            8496: bcd <= 16'h8496;
            8497: bcd <= 16'h8497;
            8498: bcd <= 16'h8498;
            8499: bcd <= 16'h8499;
            8500: bcd <= 16'h8500;
            8501: bcd <= 16'h8501;
            8502: bcd <= 16'h8502;
            8503: bcd <= 16'h8503;
            8504: bcd <= 16'h8504;
            8505: bcd <= 16'h8505;
            8506: bcd <= 16'h8506;
            8507: bcd <= 16'h8507;
            8508: bcd <= 16'h8508;
            8509: bcd <= 16'h8509;
            8510: bcd <= 16'h8510;
            8511: bcd <= 16'h8511;
            8512: bcd <= 16'h8512;
            8513: bcd <= 16'h8513;
            8514: bcd <= 16'h8514;
            8515: bcd <= 16'h8515;
            8516: bcd <= 16'h8516;
            8517: bcd <= 16'h8517;
            8518: bcd <= 16'h8518;
            8519: bcd <= 16'h8519;
            8520: bcd <= 16'h8520;
            8521: bcd <= 16'h8521;
            8522: bcd <= 16'h8522;
            8523: bcd <= 16'h8523;
            8524: bcd <= 16'h8524;
            8525: bcd <= 16'h8525;
            8526: bcd <= 16'h8526;
            8527: bcd <= 16'h8527;
            8528: bcd <= 16'h8528;
            8529: bcd <= 16'h8529;
            8530: bcd <= 16'h8530;
            8531: bcd <= 16'h8531;
            8532: bcd <= 16'h8532;
            8533: bcd <= 16'h8533;
            8534: bcd <= 16'h8534;
            8535: bcd <= 16'h8535;
            8536: bcd <= 16'h8536;
            8537: bcd <= 16'h8537;
            8538: bcd <= 16'h8538;
            8539: bcd <= 16'h8539;
            8540: bcd <= 16'h8540;
            8541: bcd <= 16'h8541;
            8542: bcd <= 16'h8542;
            8543: bcd <= 16'h8543;
            8544: bcd <= 16'h8544;
            8545: bcd <= 16'h8545;
            8546: bcd <= 16'h8546;
            8547: bcd <= 16'h8547;
            8548: bcd <= 16'h8548;
            8549: bcd <= 16'h8549;
            8550: bcd <= 16'h8550;
            8551: bcd <= 16'h8551;
            8552: bcd <= 16'h8552;
            8553: bcd <= 16'h8553;
            8554: bcd <= 16'h8554;
            8555: bcd <= 16'h8555;
            8556: bcd <= 16'h8556;
            8557: bcd <= 16'h8557;
            8558: bcd <= 16'h8558;
            8559: bcd <= 16'h8559;
            8560: bcd <= 16'h8560;
            8561: bcd <= 16'h8561;
            8562: bcd <= 16'h8562;
            8563: bcd <= 16'h8563;
            8564: bcd <= 16'h8564;
            8565: bcd <= 16'h8565;
            8566: bcd <= 16'h8566;
            8567: bcd <= 16'h8567;
            8568: bcd <= 16'h8568;
            8569: bcd <= 16'h8569;
            8570: bcd <= 16'h8570;
            8571: bcd <= 16'h8571;
            8572: bcd <= 16'h8572;
            8573: bcd <= 16'h8573;
            8574: bcd <= 16'h8574;
            8575: bcd <= 16'h8575;
            8576: bcd <= 16'h8576;
            8577: bcd <= 16'h8577;
            8578: bcd <= 16'h8578;
            8579: bcd <= 16'h8579;
            8580: bcd <= 16'h8580;
            8581: bcd <= 16'h8581;
            8582: bcd <= 16'h8582;
            8583: bcd <= 16'h8583;
            8584: bcd <= 16'h8584;
            8585: bcd <= 16'h8585;
            8586: bcd <= 16'h8586;
            8587: bcd <= 16'h8587;
            8588: bcd <= 16'h8588;
            8589: bcd <= 16'h8589;
            8590: bcd <= 16'h8590;
            8591: bcd <= 16'h8591;
            8592: bcd <= 16'h8592;
            8593: bcd <= 16'h8593;
            8594: bcd <= 16'h8594;
            8595: bcd <= 16'h8595;
            8596: bcd <= 16'h8596;
            8597: bcd <= 16'h8597;
            8598: bcd <= 16'h8598;
            8599: bcd <= 16'h8599;
            8600: bcd <= 16'h8600;
            8601: bcd <= 16'h8601;
            8602: bcd <= 16'h8602;
            8603: bcd <= 16'h8603;
            8604: bcd <= 16'h8604;
            8605: bcd <= 16'h8605;
            8606: bcd <= 16'h8606;
            8607: bcd <= 16'h8607;
            8608: bcd <= 16'h8608;
            8609: bcd <= 16'h8609;
            8610: bcd <= 16'h8610;
            8611: bcd <= 16'h8611;
            8612: bcd <= 16'h8612;
            8613: bcd <= 16'h8613;
            8614: bcd <= 16'h8614;
            8615: bcd <= 16'h8615;
            8616: bcd <= 16'h8616;
            8617: bcd <= 16'h8617;
            8618: bcd <= 16'h8618;
            8619: bcd <= 16'h8619;
            8620: bcd <= 16'h8620;
            8621: bcd <= 16'h8621;
            8622: bcd <= 16'h8622;
            8623: bcd <= 16'h8623;
            8624: bcd <= 16'h8624;
            8625: bcd <= 16'h8625;
            8626: bcd <= 16'h8626;
            8627: bcd <= 16'h8627;
            8628: bcd <= 16'h8628;
            8629: bcd <= 16'h8629;
            8630: bcd <= 16'h8630;
            8631: bcd <= 16'h8631;
            8632: bcd <= 16'h8632;
            8633: bcd <= 16'h8633;
            8634: bcd <= 16'h8634;
            8635: bcd <= 16'h8635;
            8636: bcd <= 16'h8636;
            8637: bcd <= 16'h8637;
            8638: bcd <= 16'h8638;
            8639: bcd <= 16'h8639;
            8640: bcd <= 16'h8640;
            8641: bcd <= 16'h8641;
            8642: bcd <= 16'h8642;
            8643: bcd <= 16'h8643;
            8644: bcd <= 16'h8644;
            8645: bcd <= 16'h8645;
            8646: bcd <= 16'h8646;
            8647: bcd <= 16'h8647;
            8648: bcd <= 16'h8648;
            8649: bcd <= 16'h8649;
            8650: bcd <= 16'h8650;
            8651: bcd <= 16'h8651;
            8652: bcd <= 16'h8652;
            8653: bcd <= 16'h8653;
            8654: bcd <= 16'h8654;
            8655: bcd <= 16'h8655;
            8656: bcd <= 16'h8656;
            8657: bcd <= 16'h8657;
            8658: bcd <= 16'h8658;
            8659: bcd <= 16'h8659;
            8660: bcd <= 16'h8660;
            8661: bcd <= 16'h8661;
            8662: bcd <= 16'h8662;
            8663: bcd <= 16'h8663;
            8664: bcd <= 16'h8664;
            8665: bcd <= 16'h8665;
            8666: bcd <= 16'h8666;
            8667: bcd <= 16'h8667;
            8668: bcd <= 16'h8668;
            8669: bcd <= 16'h8669;
            8670: bcd <= 16'h8670;
            8671: bcd <= 16'h8671;
            8672: bcd <= 16'h8672;
            8673: bcd <= 16'h8673;
            8674: bcd <= 16'h8674;
            8675: bcd <= 16'h8675;
            8676: bcd <= 16'h8676;
            8677: bcd <= 16'h8677;
            8678: bcd <= 16'h8678;
            8679: bcd <= 16'h8679;
            8680: bcd <= 16'h8680;
            8681: bcd <= 16'h8681;
            8682: bcd <= 16'h8682;
            8683: bcd <= 16'h8683;
            8684: bcd <= 16'h8684;
            8685: bcd <= 16'h8685;
            8686: bcd <= 16'h8686;
            8687: bcd <= 16'h8687;
            8688: bcd <= 16'h8688;
            8689: bcd <= 16'h8689;
            8690: bcd <= 16'h8690;
            8691: bcd <= 16'h8691;
            8692: bcd <= 16'h8692;
            8693: bcd <= 16'h8693;
            8694: bcd <= 16'h8694;
            8695: bcd <= 16'h8695;
            8696: bcd <= 16'h8696;
            8697: bcd <= 16'h8697;
            8698: bcd <= 16'h8698;
            8699: bcd <= 16'h8699;
            8700: bcd <= 16'h8700;
            8701: bcd <= 16'h8701;
            8702: bcd <= 16'h8702;
            8703: bcd <= 16'h8703;
            8704: bcd <= 16'h8704;
            8705: bcd <= 16'h8705;
            8706: bcd <= 16'h8706;
            8707: bcd <= 16'h8707;
            8708: bcd <= 16'h8708;
            8709: bcd <= 16'h8709;
            8710: bcd <= 16'h8710;
            8711: bcd <= 16'h8711;
            8712: bcd <= 16'h8712;
            8713: bcd <= 16'h8713;
            8714: bcd <= 16'h8714;
            8715: bcd <= 16'h8715;
            8716: bcd <= 16'h8716;
            8717: bcd <= 16'h8717;
            8718: bcd <= 16'h8718;
            8719: bcd <= 16'h8719;
            8720: bcd <= 16'h8720;
            8721: bcd <= 16'h8721;
            8722: bcd <= 16'h8722;
            8723: bcd <= 16'h8723;
            8724: bcd <= 16'h8724;
            8725: bcd <= 16'h8725;
            8726: bcd <= 16'h8726;
            8727: bcd <= 16'h8727;
            8728: bcd <= 16'h8728;
            8729: bcd <= 16'h8729;
            8730: bcd <= 16'h8730;
            8731: bcd <= 16'h8731;
            8732: bcd <= 16'h8732;
            8733: bcd <= 16'h8733;
            8734: bcd <= 16'h8734;
            8735: bcd <= 16'h8735;
            8736: bcd <= 16'h8736;
            8737: bcd <= 16'h8737;
            8738: bcd <= 16'h8738;
            8739: bcd <= 16'h8739;
            8740: bcd <= 16'h8740;
            8741: bcd <= 16'h8741;
            8742: bcd <= 16'h8742;
            8743: bcd <= 16'h8743;
            8744: bcd <= 16'h8744;
            8745: bcd <= 16'h8745;
            8746: bcd <= 16'h8746;
            8747: bcd <= 16'h8747;
            8748: bcd <= 16'h8748;
            8749: bcd <= 16'h8749;
            8750: bcd <= 16'h8750;
            8751: bcd <= 16'h8751;
            8752: bcd <= 16'h8752;
            8753: bcd <= 16'h8753;
            8754: bcd <= 16'h8754;
            8755: bcd <= 16'h8755;
            8756: bcd <= 16'h8756;
            8757: bcd <= 16'h8757;
            8758: bcd <= 16'h8758;
            8759: bcd <= 16'h8759;
            8760: bcd <= 16'h8760;
            8761: bcd <= 16'h8761;
            8762: bcd <= 16'h8762;
            8763: bcd <= 16'h8763;
            8764: bcd <= 16'h8764;
            8765: bcd <= 16'h8765;
            8766: bcd <= 16'h8766;
            8767: bcd <= 16'h8767;
            8768: bcd <= 16'h8768;
            8769: bcd <= 16'h8769;
            8770: bcd <= 16'h8770;
            8771: bcd <= 16'h8771;
            8772: bcd <= 16'h8772;
            8773: bcd <= 16'h8773;
            8774: bcd <= 16'h8774;
            8775: bcd <= 16'h8775;
            8776: bcd <= 16'h8776;
            8777: bcd <= 16'h8777;
            8778: bcd <= 16'h8778;
            8779: bcd <= 16'h8779;
            8780: bcd <= 16'h8780;
            8781: bcd <= 16'h8781;
            8782: bcd <= 16'h8782;
            8783: bcd <= 16'h8783;
            8784: bcd <= 16'h8784;
            8785: bcd <= 16'h8785;
            8786: bcd <= 16'h8786;
            8787: bcd <= 16'h8787;
            8788: bcd <= 16'h8788;
            8789: bcd <= 16'h8789;
            8790: bcd <= 16'h8790;
            8791: bcd <= 16'h8791;
            8792: bcd <= 16'h8792;
            8793: bcd <= 16'h8793;
            8794: bcd <= 16'h8794;
            8795: bcd <= 16'h8795;
            8796: bcd <= 16'h8796;
            8797: bcd <= 16'h8797;
            8798: bcd <= 16'h8798;
            8799: bcd <= 16'h8799;
            8800: bcd <= 16'h8800;
            8801: bcd <= 16'h8801;
            8802: bcd <= 16'h8802;
            8803: bcd <= 16'h8803;
            8804: bcd <= 16'h8804;
            8805: bcd <= 16'h8805;
            8806: bcd <= 16'h8806;
            8807: bcd <= 16'h8807;
            8808: bcd <= 16'h8808;
            8809: bcd <= 16'h8809;
            8810: bcd <= 16'h8810;
            8811: bcd <= 16'h8811;
            8812: bcd <= 16'h8812;
            8813: bcd <= 16'h8813;
            8814: bcd <= 16'h8814;
            8815: bcd <= 16'h8815;
            8816: bcd <= 16'h8816;
            8817: bcd <= 16'h8817;
            8818: bcd <= 16'h8818;
            8819: bcd <= 16'h8819;
            8820: bcd <= 16'h8820;
            8821: bcd <= 16'h8821;
            8822: bcd <= 16'h8822;
            8823: bcd <= 16'h8823;
            8824: bcd <= 16'h8824;
            8825: bcd <= 16'h8825;
            8826: bcd <= 16'h8826;
            8827: bcd <= 16'h8827;
            8828: bcd <= 16'h8828;
            8829: bcd <= 16'h8829;
            8830: bcd <= 16'h8830;
            8831: bcd <= 16'h8831;
            8832: bcd <= 16'h8832;
            8833: bcd <= 16'h8833;
            8834: bcd <= 16'h8834;
            8835: bcd <= 16'h8835;
            8836: bcd <= 16'h8836;
            8837: bcd <= 16'h8837;
            8838: bcd <= 16'h8838;
            8839: bcd <= 16'h8839;
            8840: bcd <= 16'h8840;
            8841: bcd <= 16'h8841;
            8842: bcd <= 16'h8842;
            8843: bcd <= 16'h8843;
            8844: bcd <= 16'h8844;
            8845: bcd <= 16'h8845;
            8846: bcd <= 16'h8846;
            8847: bcd <= 16'h8847;
            8848: bcd <= 16'h8848;
            8849: bcd <= 16'h8849;
            8850: bcd <= 16'h8850;
            8851: bcd <= 16'h8851;
            8852: bcd <= 16'h8852;
            8853: bcd <= 16'h8853;
            8854: bcd <= 16'h8854;
            8855: bcd <= 16'h8855;
            8856: bcd <= 16'h8856;
            8857: bcd <= 16'h8857;
            8858: bcd <= 16'h8858;
            8859: bcd <= 16'h8859;
            8860: bcd <= 16'h8860;
            8861: bcd <= 16'h8861;
            8862: bcd <= 16'h8862;
            8863: bcd <= 16'h8863;
            8864: bcd <= 16'h8864;
            8865: bcd <= 16'h8865;
            8866: bcd <= 16'h8866;
            8867: bcd <= 16'h8867;
            8868: bcd <= 16'h8868;
            8869: bcd <= 16'h8869;
            8870: bcd <= 16'h8870;
            8871: bcd <= 16'h8871;
            8872: bcd <= 16'h8872;
            8873: bcd <= 16'h8873;
            8874: bcd <= 16'h8874;
            8875: bcd <= 16'h8875;
            8876: bcd <= 16'h8876;
            8877: bcd <= 16'h8877;
            8878: bcd <= 16'h8878;
            8879: bcd <= 16'h8879;
            8880: bcd <= 16'h8880;
            8881: bcd <= 16'h8881;
            8882: bcd <= 16'h8882;
            8883: bcd <= 16'h8883;
            8884: bcd <= 16'h8884;
            8885: bcd <= 16'h8885;
            8886: bcd <= 16'h8886;
            8887: bcd <= 16'h8887;
            8888: bcd <= 16'h8888;
            8889: bcd <= 16'h8889;
            8890: bcd <= 16'h8890;
            8891: bcd <= 16'h8891;
            8892: bcd <= 16'h8892;
            8893: bcd <= 16'h8893;
            8894: bcd <= 16'h8894;
            8895: bcd <= 16'h8895;
            8896: bcd <= 16'h8896;
            8897: bcd <= 16'h8897;
            8898: bcd <= 16'h8898;
            8899: bcd <= 16'h8899;
            8900: bcd <= 16'h8900;
            8901: bcd <= 16'h8901;
            8902: bcd <= 16'h8902;
            8903: bcd <= 16'h8903;
            8904: bcd <= 16'h8904;
            8905: bcd <= 16'h8905;
            8906: bcd <= 16'h8906;
            8907: bcd <= 16'h8907;
            8908: bcd <= 16'h8908;
            8909: bcd <= 16'h8909;
            8910: bcd <= 16'h8910;
            8911: bcd <= 16'h8911;
            8912: bcd <= 16'h8912;
            8913: bcd <= 16'h8913;
            8914: bcd <= 16'h8914;
            8915: bcd <= 16'h8915;
            8916: bcd <= 16'h8916;
            8917: bcd <= 16'h8917;
            8918: bcd <= 16'h8918;
            8919: bcd <= 16'h8919;
            8920: bcd <= 16'h8920;
            8921: bcd <= 16'h8921;
            8922: bcd <= 16'h8922;
            8923: bcd <= 16'h8923;
            8924: bcd <= 16'h8924;
            8925: bcd <= 16'h8925;
            8926: bcd <= 16'h8926;
            8927: bcd <= 16'h8927;
            8928: bcd <= 16'h8928;
            8929: bcd <= 16'h8929;
            8930: bcd <= 16'h8930;
            8931: bcd <= 16'h8931;
            8932: bcd <= 16'h8932;
            8933: bcd <= 16'h8933;
            8934: bcd <= 16'h8934;
            8935: bcd <= 16'h8935;
            8936: bcd <= 16'h8936;
            8937: bcd <= 16'h8937;
            8938: bcd <= 16'h8938;
            8939: bcd <= 16'h8939;
            8940: bcd <= 16'h8940;
            8941: bcd <= 16'h8941;
            8942: bcd <= 16'h8942;
            8943: bcd <= 16'h8943;
            8944: bcd <= 16'h8944;
            8945: bcd <= 16'h8945;
            8946: bcd <= 16'h8946;
            8947: bcd <= 16'h8947;
            8948: bcd <= 16'h8948;
            8949: bcd <= 16'h8949;
            8950: bcd <= 16'h8950;
            8951: bcd <= 16'h8951;
            8952: bcd <= 16'h8952;
            8953: bcd <= 16'h8953;
            8954: bcd <= 16'h8954;
            8955: bcd <= 16'h8955;
            8956: bcd <= 16'h8956;
            8957: bcd <= 16'h8957;
            8958: bcd <= 16'h8958;
            8959: bcd <= 16'h8959;
            8960: bcd <= 16'h8960;
            8961: bcd <= 16'h8961;
            8962: bcd <= 16'h8962;
            8963: bcd <= 16'h8963;
            8964: bcd <= 16'h8964;
            8965: bcd <= 16'h8965;
            8966: bcd <= 16'h8966;
            8967: bcd <= 16'h8967;
            8968: bcd <= 16'h8968;
            8969: bcd <= 16'h8969;
            8970: bcd <= 16'h8970;
            8971: bcd <= 16'h8971;
            8972: bcd <= 16'h8972;
            8973: bcd <= 16'h8973;
            8974: bcd <= 16'h8974;
            8975: bcd <= 16'h8975;
            8976: bcd <= 16'h8976;
            8977: bcd <= 16'h8977;
            8978: bcd <= 16'h8978;
            8979: bcd <= 16'h8979;
            8980: bcd <= 16'h8980;
            8981: bcd <= 16'h8981;
            8982: bcd <= 16'h8982;
            8983: bcd <= 16'h8983;
            8984: bcd <= 16'h8984;
            8985: bcd <= 16'h8985;
            8986: bcd <= 16'h8986;
            8987: bcd <= 16'h8987;
            8988: bcd <= 16'h8988;
            8989: bcd <= 16'h8989;
            8990: bcd <= 16'h8990;
            8991: bcd <= 16'h8991;
            8992: bcd <= 16'h8992;
            8993: bcd <= 16'h8993;
            8994: bcd <= 16'h8994;
            8995: bcd <= 16'h8995;
            8996: bcd <= 16'h8996;
            8997: bcd <= 16'h8997;
            8998: bcd <= 16'h8998;
            8999: bcd <= 16'h8999;
            9000: bcd <= 16'h9000;
            9001: bcd <= 16'h9001;
            9002: bcd <= 16'h9002;
            9003: bcd <= 16'h9003;
            9004: bcd <= 16'h9004;
            9005: bcd <= 16'h9005;
            9006: bcd <= 16'h9006;
            9007: bcd <= 16'h9007;
            9008: bcd <= 16'h9008;
            9009: bcd <= 16'h9009;
            9010: bcd <= 16'h9010;
            9011: bcd <= 16'h9011;
            9012: bcd <= 16'h9012;
            9013: bcd <= 16'h9013;
            9014: bcd <= 16'h9014;
            9015: bcd <= 16'h9015;
            9016: bcd <= 16'h9016;
            9017: bcd <= 16'h9017;
            9018: bcd <= 16'h9018;
            9019: bcd <= 16'h9019;
            9020: bcd <= 16'h9020;
            9021: bcd <= 16'h9021;
            9022: bcd <= 16'h9022;
            9023: bcd <= 16'h9023;
            9024: bcd <= 16'h9024;
            9025: bcd <= 16'h9025;
            9026: bcd <= 16'h9026;
            9027: bcd <= 16'h9027;
            9028: bcd <= 16'h9028;
            9029: bcd <= 16'h9029;
            9030: bcd <= 16'h9030;
            9031: bcd <= 16'h9031;
            9032: bcd <= 16'h9032;
            9033: bcd <= 16'h9033;
            9034: bcd <= 16'h9034;
            9035: bcd <= 16'h9035;
            9036: bcd <= 16'h9036;
            9037: bcd <= 16'h9037;
            9038: bcd <= 16'h9038;
            9039: bcd <= 16'h9039;
            9040: bcd <= 16'h9040;
            9041: bcd <= 16'h9041;
            9042: bcd <= 16'h9042;
            9043: bcd <= 16'h9043;
            9044: bcd <= 16'h9044;
            9045: bcd <= 16'h9045;
            9046: bcd <= 16'h9046;
            9047: bcd <= 16'h9047;
            9048: bcd <= 16'h9048;
            9049: bcd <= 16'h9049;
            9050: bcd <= 16'h9050;
            9051: bcd <= 16'h9051;
            9052: bcd <= 16'h9052;
            9053: bcd <= 16'h9053;
            9054: bcd <= 16'h9054;
            9055: bcd <= 16'h9055;
            9056: bcd <= 16'h9056;
            9057: bcd <= 16'h9057;
            9058: bcd <= 16'h9058;
            9059: bcd <= 16'h9059;
            9060: bcd <= 16'h9060;
            9061: bcd <= 16'h9061;
            9062: bcd <= 16'h9062;
            9063: bcd <= 16'h9063;
            9064: bcd <= 16'h9064;
            9065: bcd <= 16'h9065;
            9066: bcd <= 16'h9066;
            9067: bcd <= 16'h9067;
            9068: bcd <= 16'h9068;
            9069: bcd <= 16'h9069;
            9070: bcd <= 16'h9070;
            9071: bcd <= 16'h9071;
            9072: bcd <= 16'h9072;
            9073: bcd <= 16'h9073;
            9074: bcd <= 16'h9074;
            9075: bcd <= 16'h9075;
            9076: bcd <= 16'h9076;
            9077: bcd <= 16'h9077;
            9078: bcd <= 16'h9078;
            9079: bcd <= 16'h9079;
            9080: bcd <= 16'h9080;
            9081: bcd <= 16'h9081;
            9082: bcd <= 16'h9082;
            9083: bcd <= 16'h9083;
            9084: bcd <= 16'h9084;
            9085: bcd <= 16'h9085;
            9086: bcd <= 16'h9086;
            9087: bcd <= 16'h9087;
            9088: bcd <= 16'h9088;
            9089: bcd <= 16'h9089;
            9090: bcd <= 16'h9090;
            9091: bcd <= 16'h9091;
            9092: bcd <= 16'h9092;
            9093: bcd <= 16'h9093;
            9094: bcd <= 16'h9094;
            9095: bcd <= 16'h9095;
            9096: bcd <= 16'h9096;
            9097: bcd <= 16'h9097;
            9098: bcd <= 16'h9098;
            9099: bcd <= 16'h9099;
            9100: bcd <= 16'h9100;
            9101: bcd <= 16'h9101;
            9102: bcd <= 16'h9102;
            9103: bcd <= 16'h9103;
            9104: bcd <= 16'h9104;
            9105: bcd <= 16'h9105;
            9106: bcd <= 16'h9106;
            9107: bcd <= 16'h9107;
            9108: bcd <= 16'h9108;
            9109: bcd <= 16'h9109;
            9110: bcd <= 16'h9110;
            9111: bcd <= 16'h9111;
            9112: bcd <= 16'h9112;
            9113: bcd <= 16'h9113;
            9114: bcd <= 16'h9114;
            9115: bcd <= 16'h9115;
            9116: bcd <= 16'h9116;
            9117: bcd <= 16'h9117;
            9118: bcd <= 16'h9118;
            9119: bcd <= 16'h9119;
            9120: bcd <= 16'h9120;
            9121: bcd <= 16'h9121;
            9122: bcd <= 16'h9122;
            9123: bcd <= 16'h9123;
            9124: bcd <= 16'h9124;
            9125: bcd <= 16'h9125;
            9126: bcd <= 16'h9126;
            9127: bcd <= 16'h9127;
            9128: bcd <= 16'h9128;
            9129: bcd <= 16'h9129;
            9130: bcd <= 16'h9130;
            9131: bcd <= 16'h9131;
            9132: bcd <= 16'h9132;
            9133: bcd <= 16'h9133;
            9134: bcd <= 16'h9134;
            9135: bcd <= 16'h9135;
            9136: bcd <= 16'h9136;
            9137: bcd <= 16'h9137;
            9138: bcd <= 16'h9138;
            9139: bcd <= 16'h9139;
            9140: bcd <= 16'h9140;
            9141: bcd <= 16'h9141;
            9142: bcd <= 16'h9142;
            9143: bcd <= 16'h9143;
            9144: bcd <= 16'h9144;
            9145: bcd <= 16'h9145;
            9146: bcd <= 16'h9146;
            9147: bcd <= 16'h9147;
            9148: bcd <= 16'h9148;
            9149: bcd <= 16'h9149;
            9150: bcd <= 16'h9150;
            9151: bcd <= 16'h9151;
            9152: bcd <= 16'h9152;
            9153: bcd <= 16'h9153;
            9154: bcd <= 16'h9154;
            9155: bcd <= 16'h9155;
            9156: bcd <= 16'h9156;
            9157: bcd <= 16'h9157;
            9158: bcd <= 16'h9158;
            9159: bcd <= 16'h9159;
            9160: bcd <= 16'h9160;
            9161: bcd <= 16'h9161;
            9162: bcd <= 16'h9162;
            9163: bcd <= 16'h9163;
            9164: bcd <= 16'h9164;
            9165: bcd <= 16'h9165;
            9166: bcd <= 16'h9166;
            9167: bcd <= 16'h9167;
            9168: bcd <= 16'h9168;
            9169: bcd <= 16'h9169;
            9170: bcd <= 16'h9170;
            9171: bcd <= 16'h9171;
            9172: bcd <= 16'h9172;
            9173: bcd <= 16'h9173;
            9174: bcd <= 16'h9174;
            9175: bcd <= 16'h9175;
            9176: bcd <= 16'h9176;
            9177: bcd <= 16'h9177;
            9178: bcd <= 16'h9178;
            9179: bcd <= 16'h9179;
            9180: bcd <= 16'h9180;
            9181: bcd <= 16'h9181;
            9182: bcd <= 16'h9182;
            9183: bcd <= 16'h9183;
            9184: bcd <= 16'h9184;
            9185: bcd <= 16'h9185;
            9186: bcd <= 16'h9186;
            9187: bcd <= 16'h9187;
            9188: bcd <= 16'h9188;
            9189: bcd <= 16'h9189;
            9190: bcd <= 16'h9190;
            9191: bcd <= 16'h9191;
            9192: bcd <= 16'h9192;
            9193: bcd <= 16'h9193;
            9194: bcd <= 16'h9194;
            9195: bcd <= 16'h9195;
            9196: bcd <= 16'h9196;
            9197: bcd <= 16'h9197;
            9198: bcd <= 16'h9198;
            9199: bcd <= 16'h9199;
            9200: bcd <= 16'h9200;
            9201: bcd <= 16'h9201;
            9202: bcd <= 16'h9202;
            9203: bcd <= 16'h9203;
            9204: bcd <= 16'h9204;
            9205: bcd <= 16'h9205;
            9206: bcd <= 16'h9206;
            9207: bcd <= 16'h9207;
            9208: bcd <= 16'h9208;
            9209: bcd <= 16'h9209;
            9210: bcd <= 16'h9210;
            9211: bcd <= 16'h9211;
            9212: bcd <= 16'h9212;
            9213: bcd <= 16'h9213;
            9214: bcd <= 16'h9214;
            9215: bcd <= 16'h9215;
            9216: bcd <= 16'h9216;
            9217: bcd <= 16'h9217;
            9218: bcd <= 16'h9218;
            9219: bcd <= 16'h9219;
            9220: bcd <= 16'h9220;
            9221: bcd <= 16'h9221;
            9222: bcd <= 16'h9222;
            9223: bcd <= 16'h9223;
            9224: bcd <= 16'h9224;
            9225: bcd <= 16'h9225;
            9226: bcd <= 16'h9226;
            9227: bcd <= 16'h9227;
            9228: bcd <= 16'h9228;
            9229: bcd <= 16'h9229;
            9230: bcd <= 16'h9230;
            9231: bcd <= 16'h9231;
            9232: bcd <= 16'h9232;
            9233: bcd <= 16'h9233;
            9234: bcd <= 16'h9234;
            9235: bcd <= 16'h9235;
            9236: bcd <= 16'h9236;
            9237: bcd <= 16'h9237;
            9238: bcd <= 16'h9238;
            9239: bcd <= 16'h9239;
            9240: bcd <= 16'h9240;
            9241: bcd <= 16'h9241;
            9242: bcd <= 16'h9242;
            9243: bcd <= 16'h9243;
            9244: bcd <= 16'h9244;
            9245: bcd <= 16'h9245;
            9246: bcd <= 16'h9246;
            9247: bcd <= 16'h9247;
            9248: bcd <= 16'h9248;
            9249: bcd <= 16'h9249;
            9250: bcd <= 16'h9250;
            9251: bcd <= 16'h9251;
            9252: bcd <= 16'h9252;
            9253: bcd <= 16'h9253;
            9254: bcd <= 16'h9254;
            9255: bcd <= 16'h9255;
            9256: bcd <= 16'h9256;
            9257: bcd <= 16'h9257;
            9258: bcd <= 16'h9258;
            9259: bcd <= 16'h9259;
            9260: bcd <= 16'h9260;
            9261: bcd <= 16'h9261;
            9262: bcd <= 16'h9262;
            9263: bcd <= 16'h9263;
            9264: bcd <= 16'h9264;
            9265: bcd <= 16'h9265;
            9266: bcd <= 16'h9266;
            9267: bcd <= 16'h9267;
            9268: bcd <= 16'h9268;
            9269: bcd <= 16'h9269;
            9270: bcd <= 16'h9270;
            9271: bcd <= 16'h9271;
            9272: bcd <= 16'h9272;
            9273: bcd <= 16'h9273;
            9274: bcd <= 16'h9274;
            9275: bcd <= 16'h9275;
            9276: bcd <= 16'h9276;
            9277: bcd <= 16'h9277;
            9278: bcd <= 16'h9278;
            9279: bcd <= 16'h9279;
            9280: bcd <= 16'h9280;
            9281: bcd <= 16'h9281;
            9282: bcd <= 16'h9282;
            9283: bcd <= 16'h9283;
            9284: bcd <= 16'h9284;
            9285: bcd <= 16'h9285;
            9286: bcd <= 16'h9286;
            9287: bcd <= 16'h9287;
            9288: bcd <= 16'h9288;
            9289: bcd <= 16'h9289;
            9290: bcd <= 16'h9290;
            9291: bcd <= 16'h9291;
            9292: bcd <= 16'h9292;
            9293: bcd <= 16'h9293;
            9294: bcd <= 16'h9294;
            9295: bcd <= 16'h9295;
            9296: bcd <= 16'h9296;
            9297: bcd <= 16'h9297;
            9298: bcd <= 16'h9298;
            9299: bcd <= 16'h9299;
            9300: bcd <= 16'h9300;
            9301: bcd <= 16'h9301;
            9302: bcd <= 16'h9302;
            9303: bcd <= 16'h9303;
            9304: bcd <= 16'h9304;
            9305: bcd <= 16'h9305;
            9306: bcd <= 16'h9306;
            9307: bcd <= 16'h9307;
            9308: bcd <= 16'h9308;
            9309: bcd <= 16'h9309;
            9310: bcd <= 16'h9310;
            9311: bcd <= 16'h9311;
            9312: bcd <= 16'h9312;
            9313: bcd <= 16'h9313;
            9314: bcd <= 16'h9314;
            9315: bcd <= 16'h9315;
            9316: bcd <= 16'h9316;
            9317: bcd <= 16'h9317;
            9318: bcd <= 16'h9318;
            9319: bcd <= 16'h9319;
            9320: bcd <= 16'h9320;
            9321: bcd <= 16'h9321;
            9322: bcd <= 16'h9322;
            9323: bcd <= 16'h9323;
            9324: bcd <= 16'h9324;
            9325: bcd <= 16'h9325;
            9326: bcd <= 16'h9326;
            9327: bcd <= 16'h9327;
            9328: bcd <= 16'h9328;
            9329: bcd <= 16'h9329;
            9330: bcd <= 16'h9330;
            9331: bcd <= 16'h9331;
            9332: bcd <= 16'h9332;
            9333: bcd <= 16'h9333;
            9334: bcd <= 16'h9334;
            9335: bcd <= 16'h9335;
            9336: bcd <= 16'h9336;
            9337: bcd <= 16'h9337;
            9338: bcd <= 16'h9338;
            9339: bcd <= 16'h9339;
            9340: bcd <= 16'h9340;
            9341: bcd <= 16'h9341;
            9342: bcd <= 16'h9342;
            9343: bcd <= 16'h9343;
            9344: bcd <= 16'h9344;
            9345: bcd <= 16'h9345;
            9346: bcd <= 16'h9346;
            9347: bcd <= 16'h9347;
            9348: bcd <= 16'h9348;
            9349: bcd <= 16'h9349;
            9350: bcd <= 16'h9350;
            9351: bcd <= 16'h9351;
            9352: bcd <= 16'h9352;
            9353: bcd <= 16'h9353;
            9354: bcd <= 16'h9354;
            9355: bcd <= 16'h9355;
            9356: bcd <= 16'h9356;
            9357: bcd <= 16'h9357;
            9358: bcd <= 16'h9358;
            9359: bcd <= 16'h9359;
            9360: bcd <= 16'h9360;
            9361: bcd <= 16'h9361;
            9362: bcd <= 16'h9362;
            9363: bcd <= 16'h9363;
            9364: bcd <= 16'h9364;
            9365: bcd <= 16'h9365;
            9366: bcd <= 16'h9366;
            9367: bcd <= 16'h9367;
            9368: bcd <= 16'h9368;
            9369: bcd <= 16'h9369;
            9370: bcd <= 16'h9370;
            9371: bcd <= 16'h9371;
            9372: bcd <= 16'h9372;
            9373: bcd <= 16'h9373;
            9374: bcd <= 16'h9374;
            9375: bcd <= 16'h9375;
            9376: bcd <= 16'h9376;
            9377: bcd <= 16'h9377;
            9378: bcd <= 16'h9378;
            9379: bcd <= 16'h9379;
            9380: bcd <= 16'h9380;
            9381: bcd <= 16'h9381;
            9382: bcd <= 16'h9382;
            9383: bcd <= 16'h9383;
            9384: bcd <= 16'h9384;
            9385: bcd <= 16'h9385;
            9386: bcd <= 16'h9386;
            9387: bcd <= 16'h9387;
            9388: bcd <= 16'h9388;
            9389: bcd <= 16'h9389;
            9390: bcd <= 16'h9390;
            9391: bcd <= 16'h9391;
            9392: bcd <= 16'h9392;
            9393: bcd <= 16'h9393;
            9394: bcd <= 16'h9394;
            9395: bcd <= 16'h9395;
            9396: bcd <= 16'h9396;
            9397: bcd <= 16'h9397;
            9398: bcd <= 16'h9398;
            9399: bcd <= 16'h9399;
            9400: bcd <= 16'h9400;
            9401: bcd <= 16'h9401;
            9402: bcd <= 16'h9402;
            9403: bcd <= 16'h9403;
            9404: bcd <= 16'h9404;
            9405: bcd <= 16'h9405;
            9406: bcd <= 16'h9406;
            9407: bcd <= 16'h9407;
            9408: bcd <= 16'h9408;
            9409: bcd <= 16'h9409;
            9410: bcd <= 16'h9410;
            9411: bcd <= 16'h9411;
            9412: bcd <= 16'h9412;
            9413: bcd <= 16'h9413;
            9414: bcd <= 16'h9414;
            9415: bcd <= 16'h9415;
            9416: bcd <= 16'h9416;
            9417: bcd <= 16'h9417;
            9418: bcd <= 16'h9418;
            9419: bcd <= 16'h9419;
            9420: bcd <= 16'h9420;
            9421: bcd <= 16'h9421;
            9422: bcd <= 16'h9422;
            9423: bcd <= 16'h9423;
            9424: bcd <= 16'h9424;
            9425: bcd <= 16'h9425;
            9426: bcd <= 16'h9426;
            9427: bcd <= 16'h9427;
            9428: bcd <= 16'h9428;
            9429: bcd <= 16'h9429;
            9430: bcd <= 16'h9430;
            9431: bcd <= 16'h9431;
            9432: bcd <= 16'h9432;
            9433: bcd <= 16'h9433;
            9434: bcd <= 16'h9434;
            9435: bcd <= 16'h9435;
            9436: bcd <= 16'h9436;
            9437: bcd <= 16'h9437;
            9438: bcd <= 16'h9438;
            9439: bcd <= 16'h9439;
            9440: bcd <= 16'h9440;
            9441: bcd <= 16'h9441;
            9442: bcd <= 16'h9442;
            9443: bcd <= 16'h9443;
            9444: bcd <= 16'h9444;
            9445: bcd <= 16'h9445;
            9446: bcd <= 16'h9446;
            9447: bcd <= 16'h9447;
            9448: bcd <= 16'h9448;
            9449: bcd <= 16'h9449;
            9450: bcd <= 16'h9450;
            9451: bcd <= 16'h9451;
            9452: bcd <= 16'h9452;
            9453: bcd <= 16'h9453;
            9454: bcd <= 16'h9454;
            9455: bcd <= 16'h9455;
            9456: bcd <= 16'h9456;
            9457: bcd <= 16'h9457;
            9458: bcd <= 16'h9458;
            9459: bcd <= 16'h9459;
            9460: bcd <= 16'h9460;
            9461: bcd <= 16'h9461;
            9462: bcd <= 16'h9462;
            9463: bcd <= 16'h9463;
            9464: bcd <= 16'h9464;
            9465: bcd <= 16'h9465;
            9466: bcd <= 16'h9466;
            9467: bcd <= 16'h9467;
            9468: bcd <= 16'h9468;
            9469: bcd <= 16'h9469;
            9470: bcd <= 16'h9470;
            9471: bcd <= 16'h9471;
            9472: bcd <= 16'h9472;
            9473: bcd <= 16'h9473;
            9474: bcd <= 16'h9474;
            9475: bcd <= 16'h9475;
            9476: bcd <= 16'h9476;
            9477: bcd <= 16'h9477;
            9478: bcd <= 16'h9478;
            9479: bcd <= 16'h9479;
            9480: bcd <= 16'h9480;
            9481: bcd <= 16'h9481;
            9482: bcd <= 16'h9482;
            9483: bcd <= 16'h9483;
            9484: bcd <= 16'h9484;
            9485: bcd <= 16'h9485;
            9486: bcd <= 16'h9486;
            9487: bcd <= 16'h9487;
            9488: bcd <= 16'h9488;
            9489: bcd <= 16'h9489;
            9490: bcd <= 16'h9490;
            9491: bcd <= 16'h9491;
            9492: bcd <= 16'h9492;
            9493: bcd <= 16'h9493;
            9494: bcd <= 16'h9494;
            9495: bcd <= 16'h9495;
            9496: bcd <= 16'h9496;
            9497: bcd <= 16'h9497;
            9498: bcd <= 16'h9498;
            9499: bcd <= 16'h9499;
            9500: bcd <= 16'h9500;
            9501: bcd <= 16'h9501;
            9502: bcd <= 16'h9502;
            9503: bcd <= 16'h9503;
            9504: bcd <= 16'h9504;
            9505: bcd <= 16'h9505;
            9506: bcd <= 16'h9506;
            9507: bcd <= 16'h9507;
            9508: bcd <= 16'h9508;
            9509: bcd <= 16'h9509;
            9510: bcd <= 16'h9510;
            9511: bcd <= 16'h9511;
            9512: bcd <= 16'h9512;
            9513: bcd <= 16'h9513;
            9514: bcd <= 16'h9514;
            9515: bcd <= 16'h9515;
            9516: bcd <= 16'h9516;
            9517: bcd <= 16'h9517;
            9518: bcd <= 16'h9518;
            9519: bcd <= 16'h9519;
            9520: bcd <= 16'h9520;
            9521: bcd <= 16'h9521;
            9522: bcd <= 16'h9522;
            9523: bcd <= 16'h9523;
            9524: bcd <= 16'h9524;
            9525: bcd <= 16'h9525;
            9526: bcd <= 16'h9526;
            9527: bcd <= 16'h9527;
            9528: bcd <= 16'h9528;
            9529: bcd <= 16'h9529;
            9530: bcd <= 16'h9530;
            9531: bcd <= 16'h9531;
            9532: bcd <= 16'h9532;
            9533: bcd <= 16'h9533;
            9534: bcd <= 16'h9534;
            9535: bcd <= 16'h9535;
            9536: bcd <= 16'h9536;
            9537: bcd <= 16'h9537;
            9538: bcd <= 16'h9538;
            9539: bcd <= 16'h9539;
            9540: bcd <= 16'h9540;
            9541: bcd <= 16'h9541;
            9542: bcd <= 16'h9542;
            9543: bcd <= 16'h9543;
            9544: bcd <= 16'h9544;
            9545: bcd <= 16'h9545;
            9546: bcd <= 16'h9546;
            9547: bcd <= 16'h9547;
            9548: bcd <= 16'h9548;
            9549: bcd <= 16'h9549;
            9550: bcd <= 16'h9550;
            9551: bcd <= 16'h9551;
            9552: bcd <= 16'h9552;
            9553: bcd <= 16'h9553;
            9554: bcd <= 16'h9554;
            9555: bcd <= 16'h9555;
            9556: bcd <= 16'h9556;
            9557: bcd <= 16'h9557;
            9558: bcd <= 16'h9558;
            9559: bcd <= 16'h9559;
            9560: bcd <= 16'h9560;
            9561: bcd <= 16'h9561;
            9562: bcd <= 16'h9562;
            9563: bcd <= 16'h9563;
            9564: bcd <= 16'h9564;
            9565: bcd <= 16'h9565;
            9566: bcd <= 16'h9566;
            9567: bcd <= 16'h9567;
            9568: bcd <= 16'h9568;
            9569: bcd <= 16'h9569;
            9570: bcd <= 16'h9570;
            9571: bcd <= 16'h9571;
            9572: bcd <= 16'h9572;
            9573: bcd <= 16'h9573;
            9574: bcd <= 16'h9574;
            9575: bcd <= 16'h9575;
            9576: bcd <= 16'h9576;
            9577: bcd <= 16'h9577;
            9578: bcd <= 16'h9578;
            9579: bcd <= 16'h9579;
            9580: bcd <= 16'h9580;
            9581: bcd <= 16'h9581;
            9582: bcd <= 16'h9582;
            9583: bcd <= 16'h9583;
            9584: bcd <= 16'h9584;
            9585: bcd <= 16'h9585;
            9586: bcd <= 16'h9586;
            9587: bcd <= 16'h9587;
            9588: bcd <= 16'h9588;
            9589: bcd <= 16'h9589;
            9590: bcd <= 16'h9590;
            9591: bcd <= 16'h9591;
            9592: bcd <= 16'h9592;
            9593: bcd <= 16'h9593;
            9594: bcd <= 16'h9594;
            9595: bcd <= 16'h9595;
            9596: bcd <= 16'h9596;
            9597: bcd <= 16'h9597;
            9598: bcd <= 16'h9598;
            9599: bcd <= 16'h9599;
            9600: bcd <= 16'h9600;
            9601: bcd <= 16'h9601;
            9602: bcd <= 16'h9602;
            9603: bcd <= 16'h9603;
            9604: bcd <= 16'h9604;
            9605: bcd <= 16'h9605;
            9606: bcd <= 16'h9606;
            9607: bcd <= 16'h9607;
            9608: bcd <= 16'h9608;
            9609: bcd <= 16'h9609;
            9610: bcd <= 16'h9610;
            9611: bcd <= 16'h9611;
            9612: bcd <= 16'h9612;
            9613: bcd <= 16'h9613;
            9614: bcd <= 16'h9614;
            9615: bcd <= 16'h9615;
            9616: bcd <= 16'h9616;
            9617: bcd <= 16'h9617;
            9618: bcd <= 16'h9618;
            9619: bcd <= 16'h9619;
            9620: bcd <= 16'h9620;
            9621: bcd <= 16'h9621;
            9622: bcd <= 16'h9622;
            9623: bcd <= 16'h9623;
            9624: bcd <= 16'h9624;
            9625: bcd <= 16'h9625;
            9626: bcd <= 16'h9626;
            9627: bcd <= 16'h9627;
            9628: bcd <= 16'h9628;
            9629: bcd <= 16'h9629;
            9630: bcd <= 16'h9630;
            9631: bcd <= 16'h9631;
            9632: bcd <= 16'h9632;
            9633: bcd <= 16'h9633;
            9634: bcd <= 16'h9634;
            9635: bcd <= 16'h9635;
            9636: bcd <= 16'h9636;
            9637: bcd <= 16'h9637;
            9638: bcd <= 16'h9638;
            9639: bcd <= 16'h9639;
            9640: bcd <= 16'h9640;
            9641: bcd <= 16'h9641;
            9642: bcd <= 16'h9642;
            9643: bcd <= 16'h9643;
            9644: bcd <= 16'h9644;
            9645: bcd <= 16'h9645;
            9646: bcd <= 16'h9646;
            9647: bcd <= 16'h9647;
            9648: bcd <= 16'h9648;
            9649: bcd <= 16'h9649;
            9650: bcd <= 16'h9650;
            9651: bcd <= 16'h9651;
            9652: bcd <= 16'h9652;
            9653: bcd <= 16'h9653;
            9654: bcd <= 16'h9654;
            9655: bcd <= 16'h9655;
            9656: bcd <= 16'h9656;
            9657: bcd <= 16'h9657;
            9658: bcd <= 16'h9658;
            9659: bcd <= 16'h9659;
            9660: bcd <= 16'h9660;
            9661: bcd <= 16'h9661;
            9662: bcd <= 16'h9662;
            9663: bcd <= 16'h9663;
            9664: bcd <= 16'h9664;
            9665: bcd <= 16'h9665;
            9666: bcd <= 16'h9666;
            9667: bcd <= 16'h9667;
            9668: bcd <= 16'h9668;
            9669: bcd <= 16'h9669;
            9670: bcd <= 16'h9670;
            9671: bcd <= 16'h9671;
            9672: bcd <= 16'h9672;
            9673: bcd <= 16'h9673;
            9674: bcd <= 16'h9674;
            9675: bcd <= 16'h9675;
            9676: bcd <= 16'h9676;
            9677: bcd <= 16'h9677;
            9678: bcd <= 16'h9678;
            9679: bcd <= 16'h9679;
            9680: bcd <= 16'h9680;
            9681: bcd <= 16'h9681;
            9682: bcd <= 16'h9682;
            9683: bcd <= 16'h9683;
            9684: bcd <= 16'h9684;
            9685: bcd <= 16'h9685;
            9686: bcd <= 16'h9686;
            9687: bcd <= 16'h9687;
            9688: bcd <= 16'h9688;
            9689: bcd <= 16'h9689;
            9690: bcd <= 16'h9690;
            9691: bcd <= 16'h9691;
            9692: bcd <= 16'h9692;
            9693: bcd <= 16'h9693;
            9694: bcd <= 16'h9694;
            9695: bcd <= 16'h9695;
            9696: bcd <= 16'h9696;
            9697: bcd <= 16'h9697;
            9698: bcd <= 16'h9698;
            9699: bcd <= 16'h9699;
            9700: bcd <= 16'h9700;
            9701: bcd <= 16'h9701;
            9702: bcd <= 16'h9702;
            9703: bcd <= 16'h9703;
            9704: bcd <= 16'h9704;
            9705: bcd <= 16'h9705;
            9706: bcd <= 16'h9706;
            9707: bcd <= 16'h9707;
            9708: bcd <= 16'h9708;
            9709: bcd <= 16'h9709;
            9710: bcd <= 16'h9710;
            9711: bcd <= 16'h9711;
            9712: bcd <= 16'h9712;
            9713: bcd <= 16'h9713;
            9714: bcd <= 16'h9714;
            9715: bcd <= 16'h9715;
            9716: bcd <= 16'h9716;
            9717: bcd <= 16'h9717;
            9718: bcd <= 16'h9718;
            9719: bcd <= 16'h9719;
            9720: bcd <= 16'h9720;
            9721: bcd <= 16'h9721;
            9722: bcd <= 16'h9722;
            9723: bcd <= 16'h9723;
            9724: bcd <= 16'h9724;
            9725: bcd <= 16'h9725;
            9726: bcd <= 16'h9726;
            9727: bcd <= 16'h9727;
            9728: bcd <= 16'h9728;
            9729: bcd <= 16'h9729;
            9730: bcd <= 16'h9730;
            9731: bcd <= 16'h9731;
            9732: bcd <= 16'h9732;
            9733: bcd <= 16'h9733;
            9734: bcd <= 16'h9734;
            9735: bcd <= 16'h9735;
            9736: bcd <= 16'h9736;
            9737: bcd <= 16'h9737;
            9738: bcd <= 16'h9738;
            9739: bcd <= 16'h9739;
            9740: bcd <= 16'h9740;
            9741: bcd <= 16'h9741;
            9742: bcd <= 16'h9742;
            9743: bcd <= 16'h9743;
            9744: bcd <= 16'h9744;
            9745: bcd <= 16'h9745;
            9746: bcd <= 16'h9746;
            9747: bcd <= 16'h9747;
            9748: bcd <= 16'h9748;
            9749: bcd <= 16'h9749;
            9750: bcd <= 16'h9750;
            9751: bcd <= 16'h9751;
            9752: bcd <= 16'h9752;
            9753: bcd <= 16'h9753;
            9754: bcd <= 16'h9754;
            9755: bcd <= 16'h9755;
            9756: bcd <= 16'h9756;
            9757: bcd <= 16'h9757;
            9758: bcd <= 16'h9758;
            9759: bcd <= 16'h9759;
            9760: bcd <= 16'h9760;
            9761: bcd <= 16'h9761;
            9762: bcd <= 16'h9762;
            9763: bcd <= 16'h9763;
            9764: bcd <= 16'h9764;
            9765: bcd <= 16'h9765;
            9766: bcd <= 16'h9766;
            9767: bcd <= 16'h9767;
            9768: bcd <= 16'h9768;
            9769: bcd <= 16'h9769;
            9770: bcd <= 16'h9770;
            9771: bcd <= 16'h9771;
            9772: bcd <= 16'h9772;
            9773: bcd <= 16'h9773;
            9774: bcd <= 16'h9774;
            9775: bcd <= 16'h9775;
            9776: bcd <= 16'h9776;
            9777: bcd <= 16'h9777;
            9778: bcd <= 16'h9778;
            9779: bcd <= 16'h9779;
            9780: bcd <= 16'h9780;
            9781: bcd <= 16'h9781;
            9782: bcd <= 16'h9782;
            9783: bcd <= 16'h9783;
            9784: bcd <= 16'h9784;
            9785: bcd <= 16'h9785;
            9786: bcd <= 16'h9786;
            9787: bcd <= 16'h9787;
            9788: bcd <= 16'h9788;
            9789: bcd <= 16'h9789;
            9790: bcd <= 16'h9790;
            9791: bcd <= 16'h9791;
            9792: bcd <= 16'h9792;
            9793: bcd <= 16'h9793;
            9794: bcd <= 16'h9794;
            9795: bcd <= 16'h9795;
            9796: bcd <= 16'h9796;
            9797: bcd <= 16'h9797;
            9798: bcd <= 16'h9798;
            9799: bcd <= 16'h9799;
            9800: bcd <= 16'h9800;
            9801: bcd <= 16'h9801;
            9802: bcd <= 16'h9802;
            9803: bcd <= 16'h9803;
            9804: bcd <= 16'h9804;
            9805: bcd <= 16'h9805;
            9806: bcd <= 16'h9806;
            9807: bcd <= 16'h9807;
            9808: bcd <= 16'h9808;
            9809: bcd <= 16'h9809;
            9810: bcd <= 16'h9810;
            9811: bcd <= 16'h9811;
            9812: bcd <= 16'h9812;
            9813: bcd <= 16'h9813;
            9814: bcd <= 16'h9814;
            9815: bcd <= 16'h9815;
            9816: bcd <= 16'h9816;
            9817: bcd <= 16'h9817;
            9818: bcd <= 16'h9818;
            9819: bcd <= 16'h9819;
            9820: bcd <= 16'h9820;
            9821: bcd <= 16'h9821;
            9822: bcd <= 16'h9822;
            9823: bcd <= 16'h9823;
            9824: bcd <= 16'h9824;
            9825: bcd <= 16'h9825;
            9826: bcd <= 16'h9826;
            9827: bcd <= 16'h9827;
            9828: bcd <= 16'h9828;
            9829: bcd <= 16'h9829;
            9830: bcd <= 16'h9830;
            9831: bcd <= 16'h9831;
            9832: bcd <= 16'h9832;
            9833: bcd <= 16'h9833;
            9834: bcd <= 16'h9834;
            9835: bcd <= 16'h9835;
            9836: bcd <= 16'h9836;
            9837: bcd <= 16'h9837;
            9838: bcd <= 16'h9838;
            9839: bcd <= 16'h9839;
            9840: bcd <= 16'h9840;
            9841: bcd <= 16'h9841;
            9842: bcd <= 16'h9842;
            9843: bcd <= 16'h9843;
            9844: bcd <= 16'h9844;
            9845: bcd <= 16'h9845;
            9846: bcd <= 16'h9846;
            9847: bcd <= 16'h9847;
            9848: bcd <= 16'h9848;
            9849: bcd <= 16'h9849;
            9850: bcd <= 16'h9850;
            9851: bcd <= 16'h9851;
            9852: bcd <= 16'h9852;
            9853: bcd <= 16'h9853;
            9854: bcd <= 16'h9854;
            9855: bcd <= 16'h9855;
            9856: bcd <= 16'h9856;
            9857: bcd <= 16'h9857;
            9858: bcd <= 16'h9858;
            9859: bcd <= 16'h9859;
            9860: bcd <= 16'h9860;
            9861: bcd <= 16'h9861;
            9862: bcd <= 16'h9862;
            9863: bcd <= 16'h9863;
            9864: bcd <= 16'h9864;
            9865: bcd <= 16'h9865;
            9866: bcd <= 16'h9866;
            9867: bcd <= 16'h9867;
            9868: bcd <= 16'h9868;
            9869: bcd <= 16'h9869;
            9870: bcd <= 16'h9870;
            9871: bcd <= 16'h9871;
            9872: bcd <= 16'h9872;
            9873: bcd <= 16'h9873;
            9874: bcd <= 16'h9874;
            9875: bcd <= 16'h9875;
            9876: bcd <= 16'h9876;
            9877: bcd <= 16'h9877;
            9878: bcd <= 16'h9878;
            9879: bcd <= 16'h9879;
            9880: bcd <= 16'h9880;
            9881: bcd <= 16'h9881;
            9882: bcd <= 16'h9882;
            9883: bcd <= 16'h9883;
            9884: bcd <= 16'h9884;
            9885: bcd <= 16'h9885;
            9886: bcd <= 16'h9886;
            9887: bcd <= 16'h9887;
            9888: bcd <= 16'h9888;
            9889: bcd <= 16'h9889;
            9890: bcd <= 16'h9890;
            9891: bcd <= 16'h9891;
            9892: bcd <= 16'h9892;
            9893: bcd <= 16'h9893;
            9894: bcd <= 16'h9894;
            9895: bcd <= 16'h9895;
            9896: bcd <= 16'h9896;
            9897: bcd <= 16'h9897;
            9898: bcd <= 16'h9898;
            9899: bcd <= 16'h9899;
            9900: bcd <= 16'h9900;
            9901: bcd <= 16'h9901;
            9902: bcd <= 16'h9902;
            9903: bcd <= 16'h9903;
            9904: bcd <= 16'h9904;
            9905: bcd <= 16'h9905;
            9906: bcd <= 16'h9906;
            9907: bcd <= 16'h9907;
            9908: bcd <= 16'h9908;
            9909: bcd <= 16'h9909;
            9910: bcd <= 16'h9910;
            9911: bcd <= 16'h9911;
            9912: bcd <= 16'h9912;
            9913: bcd <= 16'h9913;
            9914: bcd <= 16'h9914;
            9915: bcd <= 16'h9915;
            9916: bcd <= 16'h9916;
            9917: bcd <= 16'h9917;
            9918: bcd <= 16'h9918;
            9919: bcd <= 16'h9919;
            9920: bcd <= 16'h9920;
            9921: bcd <= 16'h9921;
            9922: bcd <= 16'h9922;
            9923: bcd <= 16'h9923;
            9924: bcd <= 16'h9924;
            9925: bcd <= 16'h9925;
            9926: bcd <= 16'h9926;
            9927: bcd <= 16'h9927;
            9928: bcd <= 16'h9928;
            9929: bcd <= 16'h9929;
            9930: bcd <= 16'h9930;
            9931: bcd <= 16'h9931;
            9932: bcd <= 16'h9932;
            9933: bcd <= 16'h9933;
            9934: bcd <= 16'h9934;
            9935: bcd <= 16'h9935;
            9936: bcd <= 16'h9936;
            9937: bcd <= 16'h9937;
            9938: bcd <= 16'h9938;
            9939: bcd <= 16'h9939;
            9940: bcd <= 16'h9940;
            9941: bcd <= 16'h9941;
            9942: bcd <= 16'h9942;
            9943: bcd <= 16'h9943;
            9944: bcd <= 16'h9944;
            9945: bcd <= 16'h9945;
            9946: bcd <= 16'h9946;
            9947: bcd <= 16'h9947;
            9948: bcd <= 16'h9948;
            9949: bcd <= 16'h9949;
            9950: bcd <= 16'h9950;
            9951: bcd <= 16'h9951;
            9952: bcd <= 16'h9952;
            9953: bcd <= 16'h9953;
            9954: bcd <= 16'h9954;
            9955: bcd <= 16'h9955;
            9956: bcd <= 16'h9956;
            9957: bcd <= 16'h9957;
            9958: bcd <= 16'h9958;
            9959: bcd <= 16'h9959;
            9960: bcd <= 16'h9960;
            9961: bcd <= 16'h9961;
            9962: bcd <= 16'h9962;
            9963: bcd <= 16'h9963;
            9964: bcd <= 16'h9964;
            9965: bcd <= 16'h9965;
            9966: bcd <= 16'h9966;
            9967: bcd <= 16'h9967;
            9968: bcd <= 16'h9968;
            9969: bcd <= 16'h9969;
            9970: bcd <= 16'h9970;
            9971: bcd <= 16'h9971;
            9972: bcd <= 16'h9972;
            9973: bcd <= 16'h9973;
            9974: bcd <= 16'h9974;
            9975: bcd <= 16'h9975;
            9976: bcd <= 16'h9976;
            9977: bcd <= 16'h9977;
            9978: bcd <= 16'h9978;
            9979: bcd <= 16'h9979;
            9980: bcd <= 16'h9980;
            9981: bcd <= 16'h9981;
            9982: bcd <= 16'h9982;
            9983: bcd <= 16'h9983;
            9984: bcd <= 16'h9984;
            9985: bcd <= 16'h9985;
            9986: bcd <= 16'h9986;
            9987: bcd <= 16'h9987;
            9988: bcd <= 16'h9988;
            9989: bcd <= 16'h9989;
            9990: bcd <= 16'h9990;
            9991: bcd <= 16'h9991;
            9992: bcd <= 16'h9992;
            9993: bcd <= 16'h9993;
            9994: bcd <= 16'h9994;
            9995: bcd <= 16'h9995;
            9996: bcd <= 16'h9996;
            9997: bcd <= 16'h9997;
            9998: bcd <= 16'h9998;
            9999: bcd <= 16'h9999;
            default: bcd <= 16'h0000;
        endcase
    end
endmodule 